module fft1024_core(input clk,
  input reset,
  input next,
  input [63:0] i0,
  input [63:0] i1,
  output next_out,
  output [63:0] o0,
  output [63:0] o1);

  wire [31:0] s1;
  wire [31:0] s2;
  reg s4 [19:0];
  wire s3;
  wire [63:0] s5;
  wire [31:0] s6;
  reg [63:0] s8 [15:0]; // synthesis attribute ram_style of s8 is block
  reg [63:0] s7;
  reg [63:0] s9;
  reg [31:0] s10;
  reg [31:0] s11;
  reg s13 [14:0];
  wire s12;
  reg [31:0] s14;
  reg [31:0] s15;
  reg [63:0] s17 [15:0]; // synthesis attribute ram_style of s17 is block
  reg [63:0] s16;
  reg [31:0] s18;
  reg [31:0] s19;
  wire [8:0] s20;
  wire [31:0] s21;
  reg s23 [29:0];
  wire s22;
  reg [63:0] s25 [7:0]; // synthesis attribute ram_style of s25 is block
  reg [63:0] s24;
  reg [31:0] s26;
  reg [63:0] s27;
  wire [63:0] s28;
  wire [63:0] s29;
  wire [31:0] s30;
  wire [31:0] s31;
  wire [7:0] s32;
  wire [63:0] s33;
  wire [63:0] s34;
  wire [31:0] s35;
  wire [31:0] s36;
  wire [31:0] s37;
  wire [8:0] s38;
  reg [8:0] s40 [594:0];
  wire [8:0] s39;
  reg [31:0] s41;
  reg [31:0] s42;
  wire [31:0] s43;
  wire [31:0] s44;
  reg [31:0] s45;
  reg [31:0] s46;
  reg [31:0] s47;
  reg s49 [136:0];
  wire s48;
  wire [63:0] s50;
  wire [63:0] s51;
  reg [31:0] s52;
  reg [63:0] s54 [511:0]; // synthesis attribute ram_style of s54 is block
  reg [63:0] s53;
  reg [4:0] s55;
  reg [31:0] s57 [3:0];
  wire [31:0] s56;
  reg [31:0] s59 [3:0];
  wire [31:0] s58;
  wire [63:0] s60;
  reg [31:0] s61;
  reg [31:0] s62;
  wire [31:0] s63;
  wire [31:0] s64;
  wire [6:0] s65;
  reg [31:0] s66;
  reg [31:0] s67;
  wire [63:0] s68;
  reg [31:0] s69;
  wire [31:0] s70;
  reg [3:0] s72 [10:0];
  wire [3:0] s71;
  wire [31:0] s73;
  reg [3:0] s75 [6:0];
  wire [3:0] s74;
  reg [7:0] s77 [130:0];
  wire [7:0] s76;
  reg [31:0] s78;
  wire [31:0] s79;
  wire [63:0] s80;
  wire [63:0] s81;
  reg [31:0] s82;
  reg s84 [3:0];
  wire s83;
  wire [8:0] s85;
  wire [8:0] s86;
  wire [31:0] s87;
  reg s89 [3:0];
  wire s88;
  reg [31:0] s90;
  reg [31:0] s92 [3:0];
  wire [31:0] s91;
  reg [31:0] s94 [3:0];
  wire [31:0] s93;
  wire [31:0] s95;
  wire [31:0] s96;
  wire [1:0] s97;
  wire [2:0] s98;
  wire [3:0] s99;
  wire [4:0] s100;
  wire [5:0] s101;
  wire [6:0] s102;
  wire [7:0] s103;
  reg [31:0] s104;
  wire [3:0] s105;
  reg [63:0] s106;
  reg [8:0] s107;
  wire [31:0] s108;
  wire [31:0] s109;
  reg [31:0] s110;
  wire [31:0] s111;
  wire [4:0] s112;
  reg [31:0] s113;
  reg [31:0] s114;
  reg [31:0] s116 [2:0];
  wire [31:0] s115;
  reg [31:0] s118 [2:0];
  wire [31:0] s117;
  reg [31:0] s119;
  reg [31:0] s120;
  wire [31:0] s121;
  wire [63:0] s122;
  wire [31:0] s123;
  wire [31:0] s124;
  reg [31:0] s126 [2:0];
  wire [31:0] s125;
  reg [31:0] s128 [2:0];
  wire [31:0] s127;
  reg [31:0] s129;
  reg [31:0] s130;
  wire [31:0] s131;
  reg [31:0] s132;
  reg [31:0] s133;
  reg [31:0] s135 [2:0];
  wire [31:0] s134;
  reg [31:0] s137 [2:0];
  wire [31:0] s136;
  wire [8:0] s138;
  wire [31:0] s139;
  reg [31:0] s140;
  wire [31:0] s141;
  wire [31:0] s142;
  reg [31:0] s143;
  reg [31:0] s144;
  wire [63:0] s145;
  reg [31:0] s146;
  reg [8:0] s148 [8:0];
  wire [8:0] s147;
  wire [31:0] s149;
  wire [31:0] s150;
  wire [31:0] s151;
  wire [31:0] s152;
  reg [31:0] s153;
  reg [2:0] s154;
  reg s156 [72:0];
  wire s155;
  reg [63:0] s158 [7:0]; // synthesis attribute ram_style of s158 is block
  reg [63:0] s157;
  wire [31:0] s159;
  wire [31:0] s160;
  reg [31:0] s161;
  reg [31:0] s162;
  wire [8:0] s163;
  reg [31:0] s164;
  reg [31:0] s165;
  wire [63:0] s166;
  wire [63:0] s167;
  wire [31:0] s168;
  wire [31:0] s169;
  wire [63:0] s170;
  wire [63:0] s171;
  wire [63:0] s172;
  wire [31:0] s173;
  wire [31:0] s174;
  reg [31:0] s175;
  reg s176;
  wire [31:0] s177;
  wire [31:0] s178;
  wire [31:0] s179;
  reg [31:0] s180;
  reg [31:0] s181;
  wire [31:0] s182;
  wire [31:0] s183;
  wire [63:0] s184;
  wire [63:0] s185;
  reg [1:0] s186;
  wire [3:0] s187;
  wire [1:0] s188;
  reg [31:0] s189;
  reg [8:0] s190;
  reg [4:0] s192 [269:0];
  wire [4:0] s191;
  wire [5:0] s193;
  reg [63:0] s194;
  reg [63:0] s196 [511:0]; // synthesis attribute ram_style of s196 is block
  reg [63:0] s195;
  wire [31:0] s197;
  wire [63:0] s198;
  wire [63:0] s199;
  wire [31:0] s200;
  wire [31:0] s201;
  wire [4:0] s202;
  reg [63:0] s204 [63:0]; // synthesis attribute ram_style of s204 is block
  reg [63:0] s203;
  reg [63:0] s205;
  reg s207 [67:0];
  wire s206;
  reg [31:0] s208;
  reg [31:0] s209;
  reg [31:0] s210;
  wire [31:0] s211;
  reg [31:0] s213 [3:0];
  wire [31:0] s212;
  reg [31:0] s215 [3:0];
  wire [31:0] s214;
  wire [31:0] s216;
  wire [63:0] s217;
  wire [63:0] s218;
  wire [7:0] s219;
  reg [31:0] s220;
  reg [8:0] s222 [254:0];
  wire [8:0] s221;
  reg [31:0] s223;
  wire [4:0] s224;
  reg [31:0] s226 [2:0];
  wire [31:0] s225;
  reg [31:0] s228 [2:0];
  wire [31:0] s227;
  wire [31:0] s229;
  reg [31:0] s230;
  reg [31:0] s231;
  reg [31:0] s232;
  wire [31:0] s233;
  wire [31:0] s234;
  reg [6:0] s235;
  reg [7:0] s237 [126:0];
  wire [7:0] s236;
  wire [31:0] s238;
  reg [8:0] s239;
  reg s241 [5:0];
  wire s240;
  reg [31:0] s242;
  wire [4:0] s243;
  wire [31:0] s244;
  reg [31:0] s245;
  reg [3:0] s247 [295:0];
  wire [3:0] s246;
  wire [31:0] s248;
  wire [31:0] s249;
  reg [4:0] s251 [14:0];
  wire [4:0] s250;
  reg s253 [575:0];
  wire s252;
  reg [6:0] s254;
  reg [8:0] s255;
  reg [31:0] s256;
  reg [4:0] s258 [18:0];
  wire [4:0] s257;
  wire [1:0] s259;
  wire [8:0] s260;
  reg [31:0] s261;
  reg [31:0] s262;
  reg [31:0] s263;
  wire [31:0] s264;
  wire [31:0] s265;
  wire [31:0] s266;
  reg [63:0] s268 [31:0]; // synthesis attribute ram_style of s268 is block
  reg [63:0] s267;
  reg [8:0] s269;
  wire [31:0] s270;
  wire [8:0] s271;
  reg [8:0] s273 [254:0];
  wire [8:0] s272;
  reg [31:0] s274;
  reg [31:0] s275;
  reg [31:0] s276;
  reg [31:0] s277;
  reg [31:0] s278;
  reg [8:0] s280 [29:0];
  wire [8:0] s279;
  wire [31:0] s281;
  wire [31:0] s282;
  wire [3:0] s283;
  wire [31:0] s284;
  wire [31:0] s285;
  reg [31:0] s286;
  reg [31:0] s287;
  reg [1:0] s288;
  wire [31:0] s289;
  wire [31:0] s290;
  reg s292 [261:0];
  wire s291;
  wire [31:0] s293;
  reg [31:0] s294;
  wire [31:0] s295;
  wire [31:0] s296;
  reg [31:0] s297;
  wire [31:0] s298;
  reg [63:0] s300 [127:0]; // synthesis attribute ram_style of s300 is block
  reg [63:0] s299;
  reg [31:0] s302 [3:0];
  wire [31:0] s301;
  reg [31:0] s304 [3:0];
  wire [31:0] s303;
  reg [6:0] s306 [66:0];
  wire [6:0] s305;
  wire [31:0] s307;
  reg [63:0] s309;
  reg [63:0] s308;
  reg [3:0] s310;
  wire [31:0] s311;
  reg [63:0] s312;
  wire [31:0] s313;
  reg [63:0] s315 [63:0]; // synthesis attribute ram_style of s315 is block
  reg [63:0] s314;
  wire [4:0] s316;
  wire [5:0] s317;
  reg s319 [9:0];
  wire s318;
  reg s321 [3:0];
  wire s320;
  wire [31:0] s322;
  wire [31:0] s323;
  wire [31:0] s324;
  wire [31:0] s325;
  reg s326;
  wire [31:0] s327;
  wire [31:0] s328;
  wire [63:0] s329;
  wire [63:0] s330;
  reg [63:0] s332 [31:0]; // synthesis attribute ram_style of s332 is block
  reg [63:0] s331;
  wire [63:0] s333;
  wire [1:0] s334;
  reg [31:0] s335;
  reg [63:0] s336;
  reg [31:0] s337;
  wire [31:0] s338;
  wire [63:0] s339;
  reg s341 [565:0];
  wire s340;
  wire [31:0] s342;
  wire [31:0] s343;
  wire s344;
  wire [31:0] s345;
  reg [8:0] s347 [9:0];
  wire [8:0] s346;
  reg [8:0] s349 [254:0];
  wire [8:0] s348;
  reg [31:0] s351 [2:0];
  wire [31:0] s350;
  reg [31:0] s353 [2:0];
  wire [31:0] s352;
  wire [31:0] s354;
  wire [31:0] s355;
  reg [4:0] s356;
  reg [31:0] s357;
  wire [31:0] s358;
  wire [31:0] s359;
  wire [8:0] s360;
  reg [31:0] s361;
  wire [31:0] s362;
  wire [31:0] s363;
  wire [31:0] s364;
  wire [31:0] s365;
  reg [31:0] s366;
  reg [5:0] s368 [30:0];
  wire [5:0] s367;
  reg [3:0] s369;
  wire [31:0] s370;
  wire [31:0] s371;
  reg s372;
  wire [31:0] s373;
  reg [31:0] s374;
  reg [31:0] s375;
  reg [31:0] s376;
  reg [31:0] s378 [2:0];
  wire [31:0] s377;
  reg [31:0] s380 [2:0];
  wire [31:0] s379;
  reg [7:0] s382 [585:0];
  wire [7:0] s381;
  wire [31:0] s383;
  reg [31:0] s384;
  wire [8:0] s385;
  wire [31:0] s386;
  wire [31:0] s387;
  wire [8:0] s388;
  reg [31:0] s389;
  reg [31:0] s390;
  reg [31:0] s391;
  reg s393 [5:0];
  wire s392;
  reg [31:0] s394;
  wire [31:0] s395;
  reg [31:0] s396;
  wire [31:0] s397;
  wire [31:0] s398;
  reg [31:0] s399;
  reg [31:0] s400;
  wire [31:0] s401;
  wire [31:0] s402;
  reg s404 [255:0];
  wire s403;
  reg [31:0] s405;
  reg [1:0] s407 [9:0];
  wire [1:0] s406;
  reg [63:0] s408;
  reg [63:0] s410 [511:0]; // synthesis attribute ram_style of s410 is block
  reg [63:0] s409;
  wire [4:0] s411;
  reg [31:0] s412;
  reg [31:0] s414 [3:0];
  wire [31:0] s413;
  reg [31:0] s416 [3:0];
  wire [31:0] s415;
  reg [8:0] s417;
  reg [2:0] s418;
  reg [31:0] s419;
  reg [31:0] s420;
  reg [31:0] s421;
  wire [31:0] s422;
  wire [31:0] s423;
  reg [31:0] s424;
  wire [2:0] s425;
  wire [31:0] s426;
  reg [31:0] s427;
  wire [31:0] s428;
  reg [31:0] s429;
  wire [63:0] s430;
  wire [2:0] s431;
  reg [63:0] s433 [511:0]; // synthesis attribute ram_style of s433 is block
  reg [63:0] s432;
  reg [31:0] s434;
  reg [8:0] s436 [249:0];
  wire [8:0] s435;
  wire [31:0] s437;
  wire [6:0] s438;
  reg [31:0] s439;
  reg [1:0] s440;
  reg s442 [3:0];
  wire s441;
  reg [8:0] s443;
  reg [31:0] s444;
  reg [31:0] s445;
  reg [31:0] s446;
  wire [31:0] s447;
  wire [31:0] s448;
  wire s449;
  wire [31:0] s450;
  wire [31:0] s451;
  reg [63:0] s452;
  wire [31:0] s453;
  wire [31:0] s454;
  reg [31:0] s455;
  reg [31:0] s456;
  wire [5:0] s457;
  reg [8:0] s459 [9:0];
  wire [8:0] s458;
  reg [2:0] s461 [2:0];
  wire [2:0] s460;
  reg [63:0] s462;
  wire [31:0] s463;
  wire [7:0] s464;
  reg [31:0] s465;
  wire [63:0] s466;
  wire [63:0] s467;
  wire [31:0] s468;
  reg [31:0] s469;
  reg [31:0] s470;
  wire [7:0] s471;
  wire s472;
  wire s473;
  wire s474;
  wire s475;
  wire s476;
  wire s477;
  wire s478;
  wire s479;
  reg [31:0] s481 [5:0];
  wire [31:0] s480;
  reg [31:0] s483 [5:0];
  wire [31:0] s482;
  wire [31:0] s484;
  wire [31:0] s485;
  reg [31:0] s487 [3:0];
  wire [31:0] s486;
  reg [31:0] s489 [3:0];
  wire [31:0] s488;
  reg [31:0] s491 [2:0];
  wire [31:0] s490;
  reg [31:0] s493 [2:0];
  wire [31:0] s492;
  wire [31:0] s494;
  wire [31:0] s495;
  reg [31:0] s496;
  reg [2:0] s498 [313:0];
  wire [2:0] s497;
  reg [31:0] s499;
  reg [31:0] s500;
  wire [31:0] s501;
  wire [31:0] s502;
  reg [63:0] s504 [3:0]; // synthesis attribute ram_style of s504 is block
  reg [63:0] s503;
  reg s506 [511:0];
  wire s505;
  reg [7:0] s507;
  reg [4:0] s509 [14:0];
  wire [4:0] s508;
  reg [8:0] s510;
  wire [31:0] s511;
  wire [31:0] s512;
  reg s514 [555:0];
  wire s513;
  reg [31:0] s515;
  reg [31:0] s517 [2:0];
  wire [31:0] s516;
  reg [31:0] s519 [2:0];
  wire [31:0] s518;
  wire [31:0] s520;
  reg [8:0] s522 [9:0];
  wire [8:0] s521;
  wire [3:0] s523;
  reg [5:0] s524;
  reg [31:0] s525;
  reg [2:0] s527 [6:0];
  wire [2:0] s526;
  reg s529 [11:0];
  wire s528;
  reg [8:0] s530;
  reg [8:0] s531;
  wire [31:0] s532;
  reg [7:0] s533;
  reg [31:0] s534;
  wire [63:0] s535;
  wire [63:0] s536;
  reg s538 [3:0];
  wire s537;
  wire [2:0] s539;
  reg [63:0] s540;
  reg s542 [517:0];
  wire s541;
  reg s544 [24:0];
  wire s543;
  reg [63:0] s545;
  reg [7:0] s547 [126:0];
  wire [7:0] s546;
  reg [31:0] s548;
  reg s550 [3:0];
  wire s549;
  wire [31:0] s551;
  wire [63:0] s552;
  reg [31:0] s553;
  reg [31:0] s555 [3:0];
  wire [31:0] s554;
  reg [31:0] s557 [3:0];
  wire [31:0] s556;
  reg [31:0] s559;
  reg [31:0] s558;
  reg [31:0] s561;
  reg [31:0] s560;
  wire [31:0] s562;
  wire [31:0] s563;
  wire [31:0] s564;
  reg [8:0] s566 [254:0];
  wire [8:0] s565;
  wire [31:0] s567;
  reg [31:0] s568;
  reg [31:0] s569;
  wire [63:0] s570;
  reg [31:0] s571;
  reg [31:0] s573 [2:0];
  wire [31:0] s572;
  reg [31:0] s575 [2:0];
  wire [31:0] s574;
  reg [63:0] s576;
  wire [31:0] s577;
  wire [31:0] s578;
  wire [31:0] s579;
  wire [31:0] s580;
  reg [31:0] s581;
  wire [31:0] s582;
  wire [31:0] s583;
  wire [31:0] s584;
  wire [63:0] s585;
  reg [8:0] s587 [522:0];
  wire [8:0] s586;
  reg [31:0] s589;
  reg [31:0] s588;
  reg [31:0] s591;
  reg [31:0] s590;
  wire [31:0] s592;
  wire [31:0] s593;
  reg s595 [264:0];
  wire s594;
  reg s597 [40:0];
  wire s596;
  wire [31:0] s598;
  reg [8:0] s599;
  wire [31:0] s600;
  wire [31:0] s601;
  wire [63:0] s602;
  wire [63:0] s603;
  wire [31:0] s604;
  wire [31:0] s605;
  reg [7:0] s606;
  reg [31:0] s607;
  wire [31:0] s608;
  reg [31:0] s609;
  reg [31:0] s610;
  reg [31:0] s612 [5:0];
  wire [31:0] s611;
  reg [31:0] s614 [5:0];
  wire [31:0] s613;
  reg s616 [16:0];
  wire s615;
  reg s618 [5:0];
  wire s617;
  wire [63:0] s619;
  wire [63:0] s620;
  wire [31:0] s621;
  reg [31:0] s622;
  reg [63:0] s623;
  reg [31:0] s624;
  reg [63:0] s625;
  reg [31:0] s627 [3:0];
  wire [31:0] s626;
  reg [31:0] s629 [3:0];
  wire [31:0] s628;
  wire [31:0] s630;
  wire [31:0] s631;
  reg s633 [131:0];
  wire s632;
  wire [31:0] s634;
  reg [31:0] s635;
  reg [31:0] s636;
  reg [31:0] s637;
  wire [31:0] s638;
  wire [63:0] s639;
  wire [31:0] s640;
  wire [31:0] s641;
  reg [31:0] s642;
  wire [31:0] s643;
  reg s644;
  wire [31:0] s645;
  wire [31:0] s646;
  wire [31:0] s647;
  wire [31:0] s648;
  wire [63:0] s649;
  reg [31:0] s651 [2:0];
  wire [31:0] s650;
  reg [31:0] s653 [2:0];
  wire [31:0] s652;
  reg [63:0] s655 [255:0]; // synthesis attribute ram_style of s655 is block
  reg [63:0] s654;
  wire [7:0] s656;
  reg [31:0] s657;
  reg [31:0] s658;
  reg [31:0] s660 [2:0];
  wire [31:0] s659;
  reg [31:0] s662 [2:0];
  wire [31:0] s661;
  reg [31:0] s663;
  reg [31:0] s664;
  reg [31:0] s665;
  reg [31:0] s667 [2:0];
  wire [31:0] s666;
  reg [31:0] s669 [2:0];
  wire [31:0] s668;
  wire [31:0] s670;
  wire [31:0] s671;
  wire [3:0] s672;
  wire [31:0] s673;
  reg [31:0] s675 [2:0];
  wire [31:0] s674;
  reg [31:0] s677 [2:0];
  wire [31:0] s676;
  reg [31:0] s678;
  reg [31:0] s679;
  reg [31:0] s680;
  reg [5:0] s682 [34:0];
  wire [5:0] s681;
  reg [31:0] s683;
  reg [31:0] s684;
  reg s686 [545:0];
  wire s685;
  wire [31:0] s687;
  wire [31:0] s688;
  wire [31:0] s689;
  wire [31:0] s690;
  wire [8:0] s691;
  wire s692;
  reg [31:0] s693;
  reg [31:0] s694;
  reg [31:0] s695;
  reg [31:0] s696;
  reg [31:0] s697;
  reg [31:0] s698;
  reg [31:0] s699;
  reg [63:0] s700;
  reg [31:0] s701;
  reg s703 [524:0];
  wire s702;
  reg [31:0] s704;
  reg [31:0] s705;
  reg [31:0] s706;
  reg [31:0] s707;
  wire [63:0] s708;
  wire [63:0] s709;
  reg [31:0] s711 [3:0];
  wire [31:0] s710;
  reg [31:0] s713 [3:0];
  wire [31:0] s712;
  wire [31:0] s714;
  reg [3:0] s715;
  wire [31:0] s716;
  wire [31:0] s717;
  reg [6:0] s719 [62:0];
  wire [6:0] s718;
  wire [63:0] s720;
  reg [31:0] s722 [3:0];
  wire [31:0] s721;
  reg [31:0] s724 [3:0];
  wire [31:0] s723;
  reg [63:0] s725;
  reg s727 [535:0];
  wire s726;
  wire [3:0] s728;
  reg [63:0] s730 [511:0]; // synthesis attribute ram_style of s730 is block
  reg [63:0] s729;
  wire [31:0] s731;
  reg [31:0] s732;
  wire [31:0] s733;
  wire [31:0] s734;
  wire [31:0] s735;
  wire [31:0] s736;
  reg [6:0] s738 [62:0];
  wire [6:0] s737;
  reg [31:0] s739;
  reg [31:0] s741 [2:0];
  wire [31:0] s740;
  reg [31:0] s743 [2:0];
  wire [31:0] s742;
  reg [31:0] s744;
  reg [31:0] s745;
  reg [31:0] s746;
  reg [31:0] s747;
  wire [31:0] s748;
  wire [31:0] s749;
  reg [31:0] s750;
  reg [8:0] s752 [29:0];
  wire [8:0] s751;
  reg [31:0] s753;
  reg [31:0] s754;
  wire [31:0] s755;
  reg [63:0] s756;
  reg [31:0] s757;
  reg [31:0] s758;
  reg [31:0] s759;
  reg [1:0] s760;
  wire [31:0] s761;
  reg [3:0] s763 [6:0];
  wire [3:0] s762;
  wire [31:0] s764;
  wire [31:0] s765;
  reg [31:0] s766;
  wire [31:0] s767;
  wire [8:0] s768;
  reg [31:0] s769;
  reg [31:0] s770;
  reg [31:0] s771;
  reg [31:0] s773 [3:0];
  wire [31:0] s772;
  reg [31:0] s775 [3:0];
  wire [31:0] s774;
  wire [63:0] s776;
  wire [63:0] s777;
  wire [31:0] s778;
  wire [31:0] s779;
  wire s780;
  reg [8:0] s782 [19:0];
  wire [8:0] s781;
  reg [31:0] s784 [2:0];
  wire [31:0] s783;
  reg [31:0] s786 [2:0];
  wire [31:0] s785;
  reg [31:0] s788 [3:0];
  wire [31:0] s787;
  reg [31:0] s790 [3:0];
  wire [31:0] s789;
  wire [31:0] s791;
  wire [31:0] s792;
  wire [31:0] s793;
  wire [31:0] s794;
  wire [31:0] s795;
  reg [31:0] s796;
  reg [31:0] s797;
  wire [31:0] s798;
  reg [31:0] s799;
  reg [31:0] s800;
  reg [31:0] s801;
  reg s803 [249:0];
  wire s802;
  reg [31:0] s804;
  wire [31:0] s805;
  wire [31:0] s806;
  reg s808 [3:0];
  wire s807;
  reg [31:0] s809;
  wire [31:0] s810;
  wire [31:0] s811;
  wire [31:0] s812;
  reg s814;
  reg s813;
  wire [31:0] s815;
  wire [31:0] s816;
  wire [63:0] s817;
  reg [31:0] s819;
  reg [31:0] s818;
  reg [31:0] s821;
  reg [31:0] s820;
  reg [31:0] s823 [3:0];
  wire [31:0] s822;
  reg [31:0] s825 [3:0];
  wire [31:0] s824;
  reg [31:0] s826;
  reg [31:0] s827;
  wire [63:0] s828;
  wire [63:0] s829;
  reg [31:0] s830;
  reg [31:0] s831;
  reg [5:0] s832;
  wire [63:0] s833;
  reg [63:0] s834;
  wire [4:0] s835;
  wire [31:0] s836;
  reg [7:0] s838 [15:0];
  wire [7:0] s837;
  wire s839;
  wire [31:0] s840;
  reg [31:0] s842 [3:0];
  wire [31:0] s841;
  reg [31:0] s844 [3:0];
  wire [31:0] s843;
  reg s845;
  reg [1:0] s847 [324:0];
  wire [1:0] s846;
  wire [31:0] s848;
  wire [31:0] s849;
  reg s851 [69:0];
  wire s850;
  wire [31:0] s852;
  wire [31:0] s853;
  wire [31:0] s854;
  wire [31:0] s855;
  reg [31:0] s856;
  reg [31:0] s857;
  reg [31:0] s858;
  wire [6:0] s859;
  wire [31:0] s860;
  wire [31:0] s861;
  reg [31:0] s862;
  reg [31:0] s863;
  wire [8:0] s864;
  reg s866 [7:0];
  wire s865;
  wire [31:0] s867;
  wire [31:0] s868;
  reg [31:0] s869;
  reg s871 [35:0];
  wire s870;
  wire [31:0] s872;
  wire [31:0] s873;
  wire [31:0] s874;
  wire [3:0] s875;
  wire [31:0] s876;
  wire [31:0] s877;
  reg [31:0] s878;
  reg [31:0] s880 [2:0];
  wire [31:0] s879;
  reg [31:0] s882 [2:0];
  wire [31:0] s881;
  reg [63:0] s883;
  reg [4:0] s884;
  reg [63:0] s886 [255:0]; // synthesis attribute ram_style of s886 is block
  reg [63:0] s885;
  wire [31:0] s887;
  wire [31:0] s888;
  reg [31:0] s889;
  reg [31:0] s890;
  reg [31:0] s891;
  wire [31:0] s892;
  wire [31:0] s893;
  reg [31:0] s895 [2:0];
  wire [31:0] s894;
  reg [31:0] s897 [2:0];
  wire [31:0] s896;
  reg [31:0] s898;
  wire s899;
  reg [8:0] s901 [11:0];
  wire [8:0] s900;
  reg s903 [484:0];
  wire s902;
  wire [31:0] s904;
  wire [31:0] s905;
  reg [2:0] s907 [2:0];
  wire [2:0] s906;
  wire [31:0] s908;
  wire [31:0] s909;
  reg [31:0] s910;
  wire [63:0] s911;
  wire [63:0] s912;
  wire [63:0] s913;
  reg [63:0] s914;
  reg [5:0] s916 [227:0];
  wire [5:0] s915;
  reg s918 [860:0];
  wire s917;
  wire [31:0] s919;
  wire [31:0] s920;
  wire [31:0] s921;
  reg [5:0] s923 [30:0];
  wire [5:0] s922;
  reg [31:0] s924;
  reg [31:0] s925;
  reg [63:0] s927 [511:0]; // synthesis attribute ram_style of s927 is block
  reg [63:0] s926;
  reg s929 [523:0];
  wire s928;
  wire [31:0] s930;
  reg [6:0] s932 [153:0];
  wire [6:0] s931;
  wire [31:0] s933;
  wire [31:0] s934;
  wire [31:0] s935;
  reg [8:0] s937 [9:0];
  wire [8:0] s936;
  reg [31:0] s938;
  reg [63:0] s940 [3:0]; // synthesis attribute ram_style of s940 is block
  reg [63:0] s939;
  wire [63:0] s941;
  reg [63:0] s943 [127:0]; // synthesis attribute ram_style of s943 is block
  reg [63:0] s942;
  reg [8:0] s944;
  reg [31:0] s945;
  reg s947 [337:0];
  wire s946;
  wire [63:0] s948;
  wire [31:0] s949;
  wire [8:0] s950;
  reg [31:0] s951;
  reg [31:0] s952;
  wire [31:0] s953;
  reg [31:0] s954;
  reg [31:0] s956;
  reg [31:0] s955;
  reg [31:0] s958;
  reg [31:0] s957;
  wire [31:0] s959;
  wire [31:0] s960;
  integer i;
  assign s1 = s865 ? s30 : s35;
  assign s2 = s865 ? s31 : s36;
  assign s3 = s4 [19];
  assign s5 = {s419, s375};
  assign s6 = s543 ? s622 : s856;
  assign s12 = s13 [14];
  assign s20 = {s915, s98};
  assign s21 = s668 + s379;
  assign s22 = s23 [29];
  assign s28 = $signed(s698) * $signed(32'd759250124);
  assign s29 = $signed(s699) * $signed(32'd759250124);
  assign s30 = s106[63:32];
  assign s31 = s106[31:0];
  assign s32 = s219 ^ s381;
  assign s33 = $signed(s15) * $signed(s732);
  assign s34 = $signed(s14) * $signed(s732);
  assign s35 = s9[63:32];
  assign s36 = s9[31:0];
  assign s37 = s694 + s11;
  assign s38 = {s946, s103};
  assign s39 = s40 [594];
  assign s43 = s540[63:32];
  assign s44 = s540[31:0];
  assign s48 = s49 [136];
  assign s50 = $signed(s746) * $signed(s796);
  assign s51 = $signed(s745) * $signed(s796);
  assign s56 = s57 [3];
  assign s58 = s59 [3];
  assign s60 = {s412, s744};
  assign s63 = s623[63:32];
  assign s64 = s623[31:0];
  assign s65 = {s252, 6'd0};
  assign s68 = {s78, s515};
  assign s70 = s274 + s444;
  assign s71 = s72 [10];
  assign s73 = s18 - s390;
  assign s74 = s75 [6];
  assign s76 = s77 [130];
  assign s79 = s62 - s569;
  assign s80 = $signed(s862) * $signed(s704);
  assign s81 = $signed(s863) * $signed(s704);
  assign s83 = s84 [3];
  assign s85 = {s344, s507};
  assign s86 = s531 ^ s190;
  assign s87 = s740 - s516;
  assign s88 = s89 [3];
  assign s91 = s92 [3];
  assign s93 = s94 [3];
  assign s95 = s320 ? s710 : s721;
  assign s96 = s320 ? s712 : s723;
  assign s97 = s147[8:7];
  assign s98 = s147[8:6];
  assign s99 = s147[8:5];
  assign s100 = s147[8:4];
  assign s101 = s147[8:3];
  assign s102 = s147[8:2];
  assign s103 = s147[8:1];
  assign s105 = s875 ^ s728;
  assign s108 = s83 ? s626 : s212;
  assign s109 = s83 ? s628 : s214;
  assign s111 = s543 ? s739 : s389;
  assign s112 = s411 ^ s243;
  assign s115 = s116 [2];
  assign s117 = s118 [2];
  assign s121 = s500 + s571;
  assign s122 = {s898, s164};
  assign s123 = s194[63:32];
  assign s124 = s194[31:0];
  assign s125 = s126 [2];
  assign s127 = s128 [2];
  assign s131 = s896 + s785;
  assign s134 = s135 [2];
  assign s136 = s137 [2];
  assign s138 = {s837, s318};
  assign s139 = s615 ? s951 : s130;
  assign s141 = i0[63:32];
  assign s142 = i0[31:0];
  assign s145 = {s209, s210};
  assign s147 = s148 [8];
  assign s149 = s725[63:32];
  assign s150 = s725[31:0];
  assign s151 = s62 + s569;
  assign s152 = s594 ? s361 : s337;
  assign s155 = s156 [72];
  assign s159 = s535[61:30];
  assign s160 = s536[61:30];
  assign s163 = next ? 9'd0 : s768;
  assign s166 = {s624, s45};
  assign s167 = {s120, s242};
  assign s168 = s171[61:30];
  assign s169 = s172[61:30];
  assign s170 = {s208, s439};
  assign s171 = $signed(s14) * $signed(s110);
  assign s172 = $signed(s15) * $signed(s110);
  assign s173 = s902 ? s149 : s876;
  assign s174 = s902 ? s150 : s877;
  assign s177 = s291 ? s583 : s63;
  assign s178 = s291 ? s584 : s64;
  assign s179 = s181 - s678;
  assign s182 = s12 ? s465 : s146;
  assign s183 = s758 - s456;
  assign s184 = $signed(s161) * $signed(s766);
  assign s185 = $signed(s162) * $signed(s766);
  assign s187 = s310 + 4'd1;
  assign s188 = s259 ^ s334;
  assign s191 = s192 [269];
  assign s193 = s346[5:0];
  assign s197 = s695 + s424;
  assign s198 = $signed(s863) * $signed(s680);
  assign s199 = $signed(s862) * $signed(s680);
  assign s200 = s312[63:32];
  assign s201 = s312[31:0];
  assign s202 = s917 ? s224 : s55;
  assign s206 = s207 [67];
  assign s211 = s274 - s444;
  assign s212 = s213 [3];
  assign s214 = s215 [3];
  assign s216 = s180 + s496;
  assign s217 = $signed(s162) * $signed(s693);
  assign s218 = $signed(s161) * $signed(s693);
  assign s219 = {s850, 7'd0};
  assign s221 = s222 [254];
  assign s224 = s780 ? 5'd0 : s835;
  assign s225 = s226 [2];
  assign s227 = s228 [2];
  assign s229 = s543 ? s389 : s739;
  assign s233 = s694 - s11;
  assign s234 = s46 + s297;
  assign s236 = s237 [126];
  assign s238 = s615 ? s175 : s658;
  assign s240 = s241 [5];
  assign s243 = s458[4:0];
  assign s244 = s499 - s455;
  assign s246 = s247 [295];
  assign s248 = s205[63:32];
  assign s249 = s205[31:0];
  assign s250 = s251 [14];
  assign s252 = s253 [575];
  assign s257 = s258 [18];
  assign s259 = {s928, 1'd0};
  assign s260 = s360 ^ s85;
  assign s264 = s66 + s889;
  assign s265 = s33[61:30];
  assign s266 = s34[61:30];
  assign s270 = s894 - s783;
  assign s271 = {s846, s102};
  assign s272 = s273 [254];
  assign s279 = s280 [29];
  assign s281 = s596 ? s429 : s52;
  assign s282 = s67 + s827;
  assign s283 = reset ? 4'd0 : s523;
  assign s284 = s48 ? s278 : s26;
  assign s285 = s155 ? s607 : s384;
  assign s289 = s659 - s879;
  assign s290 = s758 + s456;
  assign s291 = s292 [261];
  assign s293 = s12 ? s910 : s232;
  assign s295 = s537 ? s56 : s822;
  assign s296 = s537 ? s58 : s824;
  assign s298 = s490 - s225;
  assign s301 = s302 [3];
  assign s303 = s304 [3];
  assign s305 = s306 [66];
  assign s307 = s615 ? s130 : s951;
  assign s311 = s695 - s424;
  assign s313 = s594 ? s337 : s361;
  assign s316 = reset ? 5'd0 : s202;
  assign s317 = {s340, 5'd0};
  assign s318 = s319 [9];
  assign s320 = s321 [3];
  assign s322 = s80[61:30];
  assign s323 = s81[61:30];
  assign s324 = s576[63:32];
  assign s325 = s576[31:0];
  assign s327 = s336[63:32];
  assign s328 = s336[31:0];
  assign s329 = $signed(s399) * $signed(s657);
  assign s330 = $signed(s400) * $signed(s657);
  assign s333 = {s701, s954};
  assign o0 = s720;
  assign s334 = s586[1:0];
  assign s338 = s403 ? s374 : s10;
  assign s339 = {s143, s144};
  assign s340 = s341 [565];
  assign s342 = s22 ? s141 : s811;
  assign s343 = s22 ? s142 : s812;
  assign s344 = s269[8];
  assign s345 = s771 + s684;
  assign s346 = s347 [9];
  assign s348 = s349 [254];
  assign s350 = s351 [2];
  assign s352 = s353 [2];
  assign s354 = s902 ? s876 : s149;
  assign s355 = s902 ? s877 : s150;
  assign s358 = s50[61:30];
  assign s359 = s51[61:30];
  assign s360 = {s372, 8'd0};
  assign s362 = s644 ? 32'd0 : s469;
  assign s363 = s644 ? 32'd0 : s470;
  assign s364 = s41 - s753;
  assign s365 = s42 - s754;
  assign s367 = s368 [30];
  assign s370 = s828[61:30];
  assign s371 = s829[61:30];
  assign s373 = s702 ? s925 : s548;
  assign s377 = s378 [2];
  assign s379 = s380 [2];
  assign s381 = s382 [585];
  assign s383 = s48 ? s26 : s278;
  assign s385 = {s497, s101};
  assign s386 = s625[63:32];
  assign s387 = s625[31:0];
  assign s388 = s39 ^ s781;
  assign s392 = s393 [5];
  assign s395 = s666 - s377;
  assign s397 = s776[61:30];
  assign s398 = s777[61:30];
  assign s401 = s845 ? s588 : s955;
  assign s402 = s845 ? s590 : s957;
  assign s403 = s404 [255];
  assign s406 = s407 [9];
  assign s411 = {s513, 4'd0};
  assign s413 = s414 [3];
  assign s415 = s416 [3];
  assign s422 = s28[61:30];
  assign s423 = s29[61:30];
  assign s425 = {s726, 2'd0};
  assign s426 = s275 - s924;
  assign s428 = s48 ? s140 : s801;
  assign s430 = {s294, s82};
  assign s431 = s425 ^ s539;
  assign s435 = s436 [249];
  assign s437 = s155 ? s366 : s826;
  assign s438 = s65 ^ s859;
  assign s441 = s442 [3];
  assign s447 = s66 - s889;
  assign s448 = s770 - s683;
  assign s449 = reset ? 1'd0 : s692;
  assign s450 = s329[61:30];
  assign s451 = s330[61:30];
  assign s453 = s541 ? s799 : s286;
  assign s454 = s541 ? s800 : s287;
  assign s457 = s317 ^ s193;
  assign s458 = s459 [9];
  assign s460 = s461 [2];
  assign s463 = s115 - s650;
  assign s464 = {s472, s479, s478, s477, s476, s475, s474, s473};
  assign s466 = $signed(s609) * $signed(s637);
  assign s467 = $signed(s610) * $signed(s637);
  assign s468 = s742 + s518;
  assign s471 = s443[7:0];
  assign s472 = s443[0];
  assign s473 = s443[7];
  assign s474 = s443[6];
  assign s475 = s443[5];
  assign s476 = s443[4];
  assign s477 = s443[3];
  assign s478 = s443[2];
  assign s479 = s443[1];
  assign s480 = s481 [5];
  assign s482 = s483 [5];
  assign s484 = s807 ? s301 : s486;
  assign s485 = s807 ? s303 : s488;
  assign s486 = s487 [3];
  assign s488 = s489 [3];
  assign s490 = s491 [2];
  assign s492 = s493 [2];
  assign s494 = s757 + s938;
  assign s495 = s594 ? s421 : s427;
  assign s497 = s498 [313];
  assign s501 = s802 ? s123 : s43;
  assign s502 = s802 ? s124 : s44;
  assign s505 = s506 [511];
  assign s508 = s509 [14];
  assign s511 = s644 ? s470 : 32'd0;
  assign s512 = s644 ? s469 : 32'd0;
  assign s513 = s514 [555];
  assign s516 = s517 [2];
  assign s518 = s519 [2];
  assign s520 = s594 ? s427 : s421;
  assign s521 = s522 [9];
  assign s523 = s917 ? s672 : s310;
  assign s526 = s527 [6];
  assign s528 = s529 [11];
  assign s532 = s155 ? s384 : s607;
  assign s535 = $signed(s400) * $signed(s69);
  assign s536 = $signed(s399) * $signed(s69);
  assign s537 = s538 [3];
  assign s539 = s900[2:0];
  assign s541 = s542 [517];
  assign s543 = s544 [24];
  assign s546 = s547 [126];
  assign s549 = s550 [3];
  assign s551 = s48 ? s801 : s140;
  assign s552 = {s830, s831};
  assign s554 = s555 [3];
  assign s556 = s557 [3];
  assign s562 = s12 ? s146 : s465;
  assign s563 = s176 ? s857 : s959;
  assign s564 = s176 ? s858 : s960;
  assign s565 = s566 [254];
  assign s567 = s403 ? s394 : s231;
  assign s570 = {s276, s129};
  assign s572 = s573 [2];
  assign s574 = s575 [2];
  assign s577 = s528 ? s748 : s630;
  assign s578 = s528 ? s749 : s631;
  assign s579 = s441 ? s413 : s91;
  assign s580 = s441 ? s415 : s93;
  assign s582 = s19 + s391;
  assign s583 = s462[63:32];
  assign s584 = s462[31:0];
  assign s585 = {s220, s759};
  assign s586 = s587 [522];
  assign s592 = s67 - s827;
  assign s593 = s702 ? s548 : s925;
  assign s594 = s595 [264];
  assign s596 = s597 [40];
  assign s598 = s46 - s297;
  assign s600 = s408[63:32];
  assign s601 = s408[31:0];
  assign s602 = $signed(s610) * $signed(s357);
  assign s603 = $signed(s609) * $signed(s357);
  assign s604 = s291 ? s63 : s583;
  assign s605 = s291 ? s64 : s584;
  assign s608 = s702 ? s642 : s869;
  assign s611 = s612 [5];
  assign s613 = s614 [5];
  assign s615 = s616 [16];
  assign s617 = s618 [5];
  assign s619 = $signed(s697) * $signed(s104);
  assign s620 = $signed(s696) * $signed(s104);
  assign s621 = s500 - s571;
  assign s626 = s627 [3];
  assign s628 = s629 [3];
  assign s630 = s914[63:32];
  assign s631 = s914[31:0];
  assign s632 = s633 [131];
  assign s634 = s155 ? s826 : s366;
  assign s638 = s664 - s335;
  assign s639 = {s679, s405};
  assign s640 = s3 ? s200 : s600;
  assign s641 = s3 ? s201 : s601;
  assign s643 = s596 ? s52 : s429;
  assign s645 = s619[61:30];
  assign s646 = s620[61:30];
  assign s647 = 32'd0 - s125;
  assign s648 = 32'd0 - s127;
  assign s649 = s813 ? s308 : s552;
  assign s650 = s651 [2];
  assign s652 = s653 [2];
  assign s656 = s326 ? s464 : s471;
  assign s659 = s660 [2];
  assign s661 = s662 [2];
  assign s666 = s667 [2];
  assign s668 = s669 [2];
  assign s670 = s756[63:32];
  assign s671 = s756[31:0];
  assign s672 = s899 ? 4'd0 : s187;
  assign s673 = s275 + s924;
  assign s674 = s675 [2];
  assign s676 = s677 [2];
  assign s681 = s682 [34];
  assign s685 = s686 [545];
  assign s687 = s12 ? s232 : s910;
  assign s688 = s217[61:30];
  assign s689 = s218[61:30];
  assign s690 = s757 - s938;
  assign s691 = {s931, s97};
  assign s692 = s505 ? s839 : s326;
  assign s702 = s703 [524];
  assign s708 = {s878, s534};
  assign s709 = {s261, s262};
  assign s710 = s711 [3];
  assign s712 = s713 [3];
  assign s714 = s702 ? s869 : s642;
  assign s716 = s206 ? s670 : s324;
  assign s717 = s206 ? s671 : s325;
  assign s718 = s719 [62];
  assign s720 = {s132, s133};
  assign s721 = s722 [3];
  assign s723 = s724 [3];
  assign s726 = s727 [535];
  assign s728 = s936[3:0];
  assign s731 = s543 ? s856 : s622;
  assign s733 = s545[63:32];
  assign s734 = s545[31:0];
  assign s735 = s602[61:30];
  assign s736 = s603[61:30];
  assign s737 = s738 [62];
  assign s740 = s741 [2];
  assign s742 = s743 [2];
  assign s748 = s883[63:32];
  assign s749 = s883[31:0];
  assign s751 = s752 [29];
  assign s755 = s596 ? s245 : s446;
  assign s761 = s572 - s134;
  assign s762 = s763 [6];
  assign s764 = s41 + s753;
  assign s765 = s42 + s754;
  assign o1 = s339;
  assign s767 = s47 + s396;
  assign s768 = s443 + 9'd1;
  assign s772 = s773 [3];
  assign s774 = s775 [3];
  assign s776 = $signed(s696) * $signed(s189);
  assign s777 = $signed(s697) * $signed(s189);
  assign s778 = s180 - s496;
  assign s779 = s661 + s881;
  assign s780 = s55 == 5'd17;
  assign s781 = s782 [19];
  assign s783 = s784 [2];
  assign s785 = s786 [2];
  assign s787 = s788 [3];
  assign s789 = s790 [3];
  assign s791 = s663 - s223;
  assign s792 = s834[63:32];
  assign s793 = s834[31:0];
  assign s794 = s184[61:30];
  assign s795 = s185[61:30];
  assign s798 = s61 - s445;
  assign s802 = s803 [249];
  assign s805 = s403 ? s10 : s374;
  assign s806 = s47 - s396;
  assign s807 = s808 [3];
  assign s810 = s181 + s678;
  assign s811 = i1[63:32];
  assign s812 = i1[31:0];
  assign s815 = s870 ? s733 : s248;
  assign s816 = s870 ? s734 : s249;
  assign s817 = {s90, s420};
  assign s822 = s823 [3];
  assign s824 = s825 [3];
  assign s828 = $signed(s635) * $signed(32'd759250124);
  assign s829 = $signed(s636) * $signed(32'd759250124);
  assign s833 = {s750, s165};
  assign s835 = s55 + 5'd1;
  assign s836 = s574 + s136;
  assign s837 = s838 [15];
  assign s839 = s326 + 1'd1;
  assign s840 = s61 + s445;
  assign s841 = s842 [3];
  assign s843 = s844 [3];
  assign s846 = s847 [324];
  assign s848 = s198[61:30];
  assign s849 = s199[61:30];
  assign s850 = s851 [69];
  assign s852 = s912[61:30];
  assign s853 = s913[61:30];
  assign s854 = s466[61:30];
  assign s855 = s467[61:30];
  assign s859 = s521[6:0];
  assign s860 = s549 ? s787 : s772;
  assign s861 = s549 ? s789 : s774;
  assign s864 = {s246, s100};
  assign s865 = s866 [7];
  assign s867 = s813 ? s818 : s558;
  assign s868 = s813 ? s820 : s560;
  assign s870 = s871 [35];
  assign s872 = s663 + s223;
  assign s873 = s632 ? s908 : s386;
  assign s874 = s632 ? s909 : s387;
  assign s875 = {s685, 3'd0};
  assign s876 = s452[63:32];
  assign s877 = s452[31:0];
  assign s879 = s880 [2];
  assign s881 = s882 [2];
  assign s887 = s499 + s455;
  assign s888 = s615 ? s658 : s175;
  assign s892 = s392 ? s327 : s792;
  assign s893 = s392 ? s328 : s793;
  assign s894 = s895 [2];
  assign s896 = s897 [2];
  assign s899 = s310 == 4'd8;
  assign s900 = s901 [11];
  assign s902 = s903 [484];
  assign s904 = s88 ? s554 : s841;
  assign s905 = s88 ? s556 : s843;
  assign s906 = s907 [2];
  assign next_out = s617;
  assign s908 = s700[63:32];
  assign s909 = s700[31:0];
  assign s911 = {s769, s119};
  assign s912 = $signed(s745) * $signed(s434);
  assign s913 = $signed(s746) * $signed(s434);
  assign s915 = s916 [227];
  assign s917 = s918 [860];
  assign s919 = s596 ? s446 : s245;
  assign s920 = s22 ? s811 : s141;
  assign s921 = s22 ? s812 : s142;
  assign s922 = s923 [30];
  assign s928 = s929 [523];
  assign s930 = s403 ? s231 : s394;
  assign s931 = s932 [153];
  assign s933 = s492 + s227;
  assign s934 = s240 ? s480 : s611;
  assign s935 = s240 ? s482 : s613;
  assign s936 = s937 [9];
  assign s941 = {s376, s665};
  assign s946 = s947 [337];
  assign s948 = {s952, s553};
  assign s949 = s117 + s652;
  assign s950 = {s191, s99};
  assign s953 = s664 + s335;
  assign s959 = s27[63:32];
  assign s960 = s27[31:0];
  always @(*)
    case(s526)
      0: s153 = 32'd0;
      1: s153 = 32'd410903206;
      2: s153 = 32'd759250124;
      3: s153 = 32'd992008094;
      4: s153 = 32'd1073741824;
      5: s153 = 32'd992008094;
      6: s153 = 32'd759250124;
      7: s153 = 32'd410903206;
    endcase
  always @(*)
    case(s435)
      0: s230 = 32'd0;
      1: s230 = 32'd6588355;
      2: s230 = 32'd13176463;
      3: s230 = 32'd19764075;
      4: s230 = 32'd26350943;
      5: s230 = 32'd32936819;
      6: s230 = 32'd39521454;
      7: s230 = 32'd46104602;
      8: s230 = 32'd52686014;
      9: s230 = 32'd59265442;
      10: s230 = 32'd65842639;
      11: s230 = 32'd72417357;
      12: s230 = 32'd78989348;
      13: s230 = 32'd85558366;
      14: s230 = 32'd92124162;
      15: s230 = 32'd98686490;
      16: s230 = 32'd105245103;
      17: s230 = 32'd111799753;
      18: s230 = 32'd118350193;
      19: s230 = 32'd124896178;
      20: s230 = 32'd131437461;
      21: s230 = 32'd137973795;
      22: s230 = 32'd144504935;
      23: s230 = 32'd151030634;
      24: s230 = 32'd157550647;
      25: s230 = 32'd164064728;
      26: s230 = 32'd170572632;
      27: s230 = 32'd177074114;
      28: s230 = 32'd183568930;
      29: s230 = 32'd190056834;
      30: s230 = 32'd196537583;
      31: s230 = 32'd203010932;
      32: s230 = 32'd209476638;
      33: s230 = 32'd215934457;
      34: s230 = 32'd222384146;
      35: s230 = 32'd228825463;
      36: s230 = 32'd235258165;
      37: s230 = 32'd241682009;
      38: s230 = 32'd248096754;
      39: s230 = 32'd254502159;
      40: s230 = 32'd260897981;
      41: s230 = 32'd267283981;
      42: s230 = 32'd273659918;
      43: s230 = 32'd280025551;
      44: s230 = 32'd286380642;
      45: s230 = 32'd292724951;
      46: s230 = 32'd299058239;
      47: s230 = 32'd305380267;
      48: s230 = 32'd311690798;
      49: s230 = 32'd317989594;
      50: s230 = 32'd324276418;
      51: s230 = 32'd330551034;
      52: s230 = 32'd336813204;
      53: s230 = 32'd343062693;
      54: s230 = 32'd349299266;
      55: s230 = 32'd355522688;
      56: s230 = 32'd361732725;
      57: s230 = 32'd367929143;
      58: s230 = 32'd374111709;
      59: s230 = 32'd380280189;
      60: s230 = 32'd386434352;
      61: s230 = 32'd392573967;
      62: s230 = 32'd398698801;
      63: s230 = 32'd404808624;
      64: s230 = 32'd410903206;
      65: s230 = 32'd416982318;
      66: s230 = 32'd423045731;
      67: s230 = 32'd429093217;
      68: s230 = 32'd435124547;
      69: s230 = 32'd441139495;
      70: s230 = 32'd447137835;
      71: s230 = 32'd453119340;
      72: s230 = 32'd459083785;
      73: s230 = 32'd465030947;
      74: s230 = 32'd470960600;
      75: s230 = 32'd476872521;
      76: s230 = 32'd482766489;
      77: s230 = 32'd488642280;
      78: s230 = 32'd494499675;
      79: s230 = 32'd500338452;
      80: s230 = 32'd506158392;
      81: s230 = 32'd511959274;
      82: s230 = 32'd517740882;
      83: s230 = 32'd523502998;
      84: s230 = 32'd529245403;
      85: s230 = 32'd534967883;
      86: s230 = 32'd540670222;
      87: s230 = 32'd546352205;
      88: s230 = 32'd552013618;
      89: s230 = 32'd557654248;
      90: s230 = 32'd563273882;
      91: s230 = 32'd568872310;
      92: s230 = 32'd574449320;
      93: s230 = 32'd580004702;
      94: s230 = 32'd585538247;
      95: s230 = 32'd591049747;
      96: s230 = 32'd596538995;
      97: s230 = 32'd602005783;
      98: s230 = 32'd607449906;
      99: s230 = 32'd612871159;
      100: s230 = 32'd618269337;
      101: s230 = 32'd623644238;
      102: s230 = 32'd628995659;
      103: s230 = 32'd634323399;
      104: s230 = 32'd639627257;
      105: s230 = 32'd644907034;
      106: s230 = 32'd650162530;
      107: s230 = 32'd655393547;
      108: s230 = 32'd660599890;
      109: s230 = 32'd665781361;
      110: s230 = 32'd670937766;
      111: s230 = 32'd676068911;
      112: s230 = 32'd681174602;
      113: s230 = 32'd686254647;
      114: s230 = 32'd691308855;
      115: s230 = 32'd696337035;
      116: s230 = 32'd701338999;
      117: s230 = 32'd706314558;
      118: s230 = 32'd711263525;
      119: s230 = 32'd716185713;
      120: s230 = 32'd721080937;
      121: s230 = 32'd725949012;
      122: s230 = 32'd730789756;
      123: s230 = 32'd735602987;
      124: s230 = 32'd740388522;
      125: s230 = 32'd745146182;
      126: s230 = 32'd749875787;
      127: s230 = 32'd754577161;
      128: s230 = 32'd759250124;
      129: s230 = 32'd763894503;
      130: s230 = 32'd768510121;
      131: s230 = 32'd773096806;
      132: s230 = 32'd777654383;
      133: s230 = 32'd782182683;
      134: s230 = 32'd786681534;
      135: s230 = 32'd791150766;
      136: s230 = 32'd795590212;
      137: s230 = 32'd799999705;
      138: s230 = 32'd804379078;
      139: s230 = 32'd808728167;
      140: s230 = 32'd813046807;
      141: s230 = 32'd817334837;
      142: s230 = 32'd821592095;
      143: s230 = 32'd825818420;
      144: s230 = 32'd830013654;
      145: s230 = 32'd834177638;
      146: s230 = 32'd838310215;
      147: s230 = 32'd842411231;
      148: s230 = 32'd846480531;
      149: s230 = 32'd850517961;
      150: s230 = 32'd854523369;
      151: s230 = 32'd858496605;
      152: s230 = 32'd862437519;
      153: s230 = 32'd866345963;
      154: s230 = 32'd870221790;
      155: s230 = 32'd874064853;
      156: s230 = 32'd877875008;
      157: s230 = 32'd881652112;
      158: s230 = 32'd885396022;
      159: s230 = 32'd889106597;
      160: s230 = 32'd892783698;
      161: s230 = 32'd896427186;
      162: s230 = 32'd900036924;
      163: s230 = 32'd903612776;
      164: s230 = 32'd907154608;
      165: s230 = 32'd910662286;
      166: s230 = 32'd914135677;
      167: s230 = 32'd917574653;
      168: s230 = 32'd920979082;
      169: s230 = 32'd924348836;
      170: s230 = 32'd927683790;
      171: s230 = 32'd930983817;
      172: s230 = 32'd934248792;
      173: s230 = 32'd937478594;
      174: s230 = 32'd940673100;
      175: s230 = 32'd943832191;
      176: s230 = 32'd946955747;
      177: s230 = 32'd950043650;
      178: s230 = 32'd953095785;
      179: s230 = 32'd956112036;
      180: s230 = 32'd959092290;
      181: s230 = 32'd962036435;
      182: s230 = 32'd964944359;
      183: s230 = 32'd967815955;
      184: s230 = 32'd970651112;
      185: s230 = 32'd973449725;
      186: s230 = 32'd976211688;
      187: s230 = 32'd978936897;
      188: s230 = 32'd981625250;
      189: s230 = 32'd984276645;
      190: s230 = 32'd986890983;
      191: s230 = 32'd989468165;
      192: s230 = 32'd992008094;
      193: s230 = 32'd994510674;
      194: s230 = 32'd996975812;
      195: s230 = 32'd999403414;
      196: s230 = 32'd1001793389;
      197: s230 = 32'd1004145647;
      198: s230 = 32'd1006460100;
      199: s230 = 32'd1008736660;
      200: s230 = 32'd1010975241;
      201: s230 = 32'd1013175760;
      202: s230 = 32'd1015338134;
      203: s230 = 32'd1017462280;
      204: s230 = 32'd1019548120;
      205: s230 = 32'd1021595574;
      206: s230 = 32'd1023604566;
      207: s230 = 32'd1025575020;
      208: s230 = 32'd1027506861;
      209: s230 = 32'd1029400017;
      210: s230 = 32'd1031254417;
      211: s230 = 32'd1033069991;
      212: s230 = 32'd1034846670;
      213: s230 = 32'd1036584388;
      214: s230 = 32'd1038283079;
      215: s230 = 32'd1039942680;
      216: s230 = 32'd1041563127;
      217: s230 = 32'd1043144359;
      218: s230 = 32'd1044686318;
      219: s230 = 32'd1046188946;
      220: s230 = 32'd1047652184;
      221: s230 = 32'd1049075979;
      222: s230 = 32'd1050460278;
      223: s230 = 32'd1051805026;
      224: s230 = 32'd1053110175;
      225: s230 = 32'd1054375675;
      226: s230 = 32'd1055601479;
      227: s230 = 32'd1056787539;
      228: s230 = 32'd1057933812;
      229: s230 = 32'd1059040255;
      230: s230 = 32'd1060106825;
      231: s230 = 32'd1061133483;
      232: s230 = 32'd1062120190;
      233: s230 = 32'd1063066908;
      234: s230 = 32'd1063973603;
      235: s230 = 32'd1064840239;
      236: s230 = 32'd1065666785;
      237: s230 = 32'd1066453209;
      238: s230 = 32'd1067199482;
      239: s230 = 32'd1067905576;
      240: s230 = 32'd1068571463;
      241: s230 = 32'd1069197119;
      242: s230 = 32'd1069782521;
      243: s230 = 32'd1070327646;
      244: s230 = 32'd1070832474;
      245: s230 = 32'd1071296985;
      246: s230 = 32'd1071721163;
      247: s230 = 32'd1072104991;
      248: s230 = 32'd1072448454;
      249: s230 = 32'd1072751541;
      250: s230 = 32'd1073014239;
      251: s230 = 32'd1073236539;
      252: s230 = 32'd1073418433;
      253: s230 = 32'd1073559912;
      254: s230 = 32'd1073660973;
      255: s230 = 32'd1073721611;
      256: s230 = 32'd1073741824;
      257: s230 = 32'd1073721611;
      258: s230 = 32'd1073660973;
      259: s230 = 32'd1073559912;
      260: s230 = 32'd1073418433;
      261: s230 = 32'd1073236539;
      262: s230 = 32'd1073014239;
      263: s230 = 32'd1072751541;
      264: s230 = 32'd1072448454;
      265: s230 = 32'd1072104991;
      266: s230 = 32'd1071721163;
      267: s230 = 32'd1071296985;
      268: s230 = 32'd1070832474;
      269: s230 = 32'd1070327646;
      270: s230 = 32'd1069782521;
      271: s230 = 32'd1069197119;
      272: s230 = 32'd1068571463;
      273: s230 = 32'd1067905576;
      274: s230 = 32'd1067199482;
      275: s230 = 32'd1066453209;
      276: s230 = 32'd1065666785;
      277: s230 = 32'd1064840239;
      278: s230 = 32'd1063973603;
      279: s230 = 32'd1063066908;
      280: s230 = 32'd1062120190;
      281: s230 = 32'd1061133483;
      282: s230 = 32'd1060106825;
      283: s230 = 32'd1059040255;
      284: s230 = 32'd1057933812;
      285: s230 = 32'd1056787539;
      286: s230 = 32'd1055601479;
      287: s230 = 32'd1054375675;
      288: s230 = 32'd1053110175;
      289: s230 = 32'd1051805026;
      290: s230 = 32'd1050460278;
      291: s230 = 32'd1049075979;
      292: s230 = 32'd1047652184;
      293: s230 = 32'd1046188946;
      294: s230 = 32'd1044686318;
      295: s230 = 32'd1043144359;
      296: s230 = 32'd1041563127;
      297: s230 = 32'd1039942680;
      298: s230 = 32'd1038283079;
      299: s230 = 32'd1036584388;
      300: s230 = 32'd1034846670;
      301: s230 = 32'd1033069991;
      302: s230 = 32'd1031254417;
      303: s230 = 32'd1029400017;
      304: s230 = 32'd1027506861;
      305: s230 = 32'd1025575020;
      306: s230 = 32'd1023604566;
      307: s230 = 32'd1021595574;
      308: s230 = 32'd1019548120;
      309: s230 = 32'd1017462280;
      310: s230 = 32'd1015338134;
      311: s230 = 32'd1013175760;
      312: s230 = 32'd1010975241;
      313: s230 = 32'd1008736660;
      314: s230 = 32'd1006460100;
      315: s230 = 32'd1004145647;
      316: s230 = 32'd1001793389;
      317: s230 = 32'd999403414;
      318: s230 = 32'd996975812;
      319: s230 = 32'd994510674;
      320: s230 = 32'd992008094;
      321: s230 = 32'd989468165;
      322: s230 = 32'd986890983;
      323: s230 = 32'd984276645;
      324: s230 = 32'd981625250;
      325: s230 = 32'd978936897;
      326: s230 = 32'd976211688;
      327: s230 = 32'd973449725;
      328: s230 = 32'd970651112;
      329: s230 = 32'd967815955;
      330: s230 = 32'd964944359;
      331: s230 = 32'd962036435;
      332: s230 = 32'd959092290;
      333: s230 = 32'd956112036;
      334: s230 = 32'd953095785;
      335: s230 = 32'd950043650;
      336: s230 = 32'd946955747;
      337: s230 = 32'd943832191;
      338: s230 = 32'd940673100;
      339: s230 = 32'd937478594;
      340: s230 = 32'd934248792;
      341: s230 = 32'd930983817;
      342: s230 = 32'd927683790;
      343: s230 = 32'd924348836;
      344: s230 = 32'd920979082;
      345: s230 = 32'd917574653;
      346: s230 = 32'd914135677;
      347: s230 = 32'd910662286;
      348: s230 = 32'd907154608;
      349: s230 = 32'd903612776;
      350: s230 = 32'd900036924;
      351: s230 = 32'd896427186;
      352: s230 = 32'd892783698;
      353: s230 = 32'd889106597;
      354: s230 = 32'd885396022;
      355: s230 = 32'd881652112;
      356: s230 = 32'd877875008;
      357: s230 = 32'd874064853;
      358: s230 = 32'd870221790;
      359: s230 = 32'd866345963;
      360: s230 = 32'd862437519;
      361: s230 = 32'd858496605;
      362: s230 = 32'd854523369;
      363: s230 = 32'd850517961;
      364: s230 = 32'd846480531;
      365: s230 = 32'd842411231;
      366: s230 = 32'd838310215;
      367: s230 = 32'd834177638;
      368: s230 = 32'd830013654;
      369: s230 = 32'd825818420;
      370: s230 = 32'd821592095;
      371: s230 = 32'd817334837;
      372: s230 = 32'd813046807;
      373: s230 = 32'd808728167;
      374: s230 = 32'd804379078;
      375: s230 = 32'd799999705;
      376: s230 = 32'd795590212;
      377: s230 = 32'd791150766;
      378: s230 = 32'd786681534;
      379: s230 = 32'd782182683;
      380: s230 = 32'd777654383;
      381: s230 = 32'd773096806;
      382: s230 = 32'd768510121;
      383: s230 = 32'd763894503;
      384: s230 = 32'd759250124;
      385: s230 = 32'd754577161;
      386: s230 = 32'd749875787;
      387: s230 = 32'd745146182;
      388: s230 = 32'd740388522;
      389: s230 = 32'd735602987;
      390: s230 = 32'd730789756;
      391: s230 = 32'd725949012;
      392: s230 = 32'd721080937;
      393: s230 = 32'd716185713;
      394: s230 = 32'd711263525;
      395: s230 = 32'd706314558;
      396: s230 = 32'd701338999;
      397: s230 = 32'd696337035;
      398: s230 = 32'd691308855;
      399: s230 = 32'd686254647;
      400: s230 = 32'd681174602;
      401: s230 = 32'd676068911;
      402: s230 = 32'd670937766;
      403: s230 = 32'd665781361;
      404: s230 = 32'd660599890;
      405: s230 = 32'd655393547;
      406: s230 = 32'd650162530;
      407: s230 = 32'd644907034;
      408: s230 = 32'd639627257;
      409: s230 = 32'd634323399;
      410: s230 = 32'd628995659;
      411: s230 = 32'd623644238;
      412: s230 = 32'd618269337;
      413: s230 = 32'd612871159;
      414: s230 = 32'd607449906;
      415: s230 = 32'd602005783;
      416: s230 = 32'd596538995;
      417: s230 = 32'd591049747;
      418: s230 = 32'd585538247;
      419: s230 = 32'd580004702;
      420: s230 = 32'd574449320;
      421: s230 = 32'd568872310;
      422: s230 = 32'd563273882;
      423: s230 = 32'd557654248;
      424: s230 = 32'd552013618;
      425: s230 = 32'd546352205;
      426: s230 = 32'd540670222;
      427: s230 = 32'd534967883;
      428: s230 = 32'd529245403;
      429: s230 = 32'd523502998;
      430: s230 = 32'd517740882;
      431: s230 = 32'd511959274;
      432: s230 = 32'd506158392;
      433: s230 = 32'd500338452;
      434: s230 = 32'd494499675;
      435: s230 = 32'd488642280;
      436: s230 = 32'd482766489;
      437: s230 = 32'd476872521;
      438: s230 = 32'd470960600;
      439: s230 = 32'd465030947;
      440: s230 = 32'd459083785;
      441: s230 = 32'd453119340;
      442: s230 = 32'd447137835;
      443: s230 = 32'd441139495;
      444: s230 = 32'd435124547;
      445: s230 = 32'd429093217;
      446: s230 = 32'd423045731;
      447: s230 = 32'd416982318;
      448: s230 = 32'd410903206;
      449: s230 = 32'd404808624;
      450: s230 = 32'd398698801;
      451: s230 = 32'd392573967;
      452: s230 = 32'd386434352;
      453: s230 = 32'd380280189;
      454: s230 = 32'd374111709;
      455: s230 = 32'd367929143;
      456: s230 = 32'd361732725;
      457: s230 = 32'd355522688;
      458: s230 = 32'd349299266;
      459: s230 = 32'd343062693;
      460: s230 = 32'd336813204;
      461: s230 = 32'd330551034;
      462: s230 = 32'd324276418;
      463: s230 = 32'd317989594;
      464: s230 = 32'd311690798;
      465: s230 = 32'd305380267;
      466: s230 = 32'd299058239;
      467: s230 = 32'd292724951;
      468: s230 = 32'd286380642;
      469: s230 = 32'd280025551;
      470: s230 = 32'd273659918;
      471: s230 = 32'd267283981;
      472: s230 = 32'd260897981;
      473: s230 = 32'd254502159;
      474: s230 = 32'd248096754;
      475: s230 = 32'd241682009;
      476: s230 = 32'd235258165;
      477: s230 = 32'd228825463;
      478: s230 = 32'd222384146;
      479: s230 = 32'd215934457;
      480: s230 = 32'd209476638;
      481: s230 = 32'd203010932;
      482: s230 = 32'd196537583;
      483: s230 = 32'd190056834;
      484: s230 = 32'd183568930;
      485: s230 = 32'd177074114;
      486: s230 = 32'd170572632;
      487: s230 = 32'd164064728;
      488: s230 = 32'd157550647;
      489: s230 = 32'd151030634;
      490: s230 = 32'd144504935;
      491: s230 = 32'd137973795;
      492: s230 = 32'd131437461;
      493: s230 = 32'd124896178;
      494: s230 = 32'd118350193;
      495: s230 = 32'd111799753;
      496: s230 = 32'd105245103;
      497: s230 = 32'd98686490;
      498: s230 = 32'd92124162;
      499: s230 = 32'd85558366;
      500: s230 = 32'd78989348;
      501: s230 = 32'd72417357;
      502: s230 = 32'd65842639;
      503: s230 = 32'd59265442;
      504: s230 = 32'd52686014;
      505: s230 = 32'd46104602;
      506: s230 = 32'd39521454;
      507: s230 = 32'd32936819;
      508: s230 = 32'd26350943;
      509: s230 = 32'd19764075;
      510: s230 = 32'd13176463;
      511: s230 = 32'd6588355;
    endcase
  always @(*)
    case(s76)
      0: s256 = 32'd0;
      1: s256 = 32'd13176463;
      2: s256 = 32'd26350943;
      3: s256 = 32'd39521454;
      4: s256 = 32'd52686014;
      5: s256 = 32'd65842639;
      6: s256 = 32'd78989348;
      7: s256 = 32'd92124162;
      8: s256 = 32'd105245103;
      9: s256 = 32'd118350193;
      10: s256 = 32'd131437461;
      11: s256 = 32'd144504935;
      12: s256 = 32'd157550647;
      13: s256 = 32'd170572632;
      14: s256 = 32'd183568930;
      15: s256 = 32'd196537583;
      16: s256 = 32'd209476638;
      17: s256 = 32'd222384146;
      18: s256 = 32'd235258165;
      19: s256 = 32'd248096754;
      20: s256 = 32'd260897981;
      21: s256 = 32'd273659918;
      22: s256 = 32'd286380642;
      23: s256 = 32'd299058239;
      24: s256 = 32'd311690798;
      25: s256 = 32'd324276418;
      26: s256 = 32'd336813204;
      27: s256 = 32'd349299266;
      28: s256 = 32'd361732725;
      29: s256 = 32'd374111709;
      30: s256 = 32'd386434352;
      31: s256 = 32'd398698801;
      32: s256 = 32'd410903206;
      33: s256 = 32'd423045731;
      34: s256 = 32'd435124547;
      35: s256 = 32'd447137835;
      36: s256 = 32'd459083785;
      37: s256 = 32'd470960600;
      38: s256 = 32'd482766489;
      39: s256 = 32'd494499675;
      40: s256 = 32'd506158392;
      41: s256 = 32'd517740882;
      42: s256 = 32'd529245403;
      43: s256 = 32'd540670222;
      44: s256 = 32'd552013618;
      45: s256 = 32'd563273882;
      46: s256 = 32'd574449320;
      47: s256 = 32'd585538247;
      48: s256 = 32'd596538995;
      49: s256 = 32'd607449906;
      50: s256 = 32'd618269337;
      51: s256 = 32'd628995659;
      52: s256 = 32'd639627257;
      53: s256 = 32'd650162530;
      54: s256 = 32'd660599890;
      55: s256 = 32'd670937766;
      56: s256 = 32'd681174602;
      57: s256 = 32'd691308855;
      58: s256 = 32'd701338999;
      59: s256 = 32'd711263525;
      60: s256 = 32'd721080937;
      61: s256 = 32'd730789756;
      62: s256 = 32'd740388522;
      63: s256 = 32'd749875787;
      64: s256 = 32'd759250124;
      65: s256 = 32'd768510121;
      66: s256 = 32'd777654383;
      67: s256 = 32'd786681534;
      68: s256 = 32'd795590212;
      69: s256 = 32'd804379078;
      70: s256 = 32'd813046807;
      71: s256 = 32'd821592095;
      72: s256 = 32'd830013654;
      73: s256 = 32'd838310215;
      74: s256 = 32'd846480531;
      75: s256 = 32'd854523369;
      76: s256 = 32'd862437519;
      77: s256 = 32'd870221790;
      78: s256 = 32'd877875008;
      79: s256 = 32'd885396022;
      80: s256 = 32'd892783698;
      81: s256 = 32'd900036924;
      82: s256 = 32'd907154608;
      83: s256 = 32'd914135677;
      84: s256 = 32'd920979082;
      85: s256 = 32'd927683790;
      86: s256 = 32'd934248792;
      87: s256 = 32'd940673100;
      88: s256 = 32'd946955747;
      89: s256 = 32'd953095785;
      90: s256 = 32'd959092290;
      91: s256 = 32'd964944359;
      92: s256 = 32'd970651112;
      93: s256 = 32'd976211688;
      94: s256 = 32'd981625250;
      95: s256 = 32'd986890983;
      96: s256 = 32'd992008094;
      97: s256 = 32'd996975812;
      98: s256 = 32'd1001793389;
      99: s256 = 32'd1006460100;
      100: s256 = 32'd1010975241;
      101: s256 = 32'd1015338134;
      102: s256 = 32'd1019548120;
      103: s256 = 32'd1023604566;
      104: s256 = 32'd1027506861;
      105: s256 = 32'd1031254417;
      106: s256 = 32'd1034846670;
      107: s256 = 32'd1038283079;
      108: s256 = 32'd1041563127;
      109: s256 = 32'd1044686318;
      110: s256 = 32'd1047652184;
      111: s256 = 32'd1050460278;
      112: s256 = 32'd1053110175;
      113: s256 = 32'd1055601479;
      114: s256 = 32'd1057933812;
      115: s256 = 32'd1060106825;
      116: s256 = 32'd1062120190;
      117: s256 = 32'd1063973603;
      118: s256 = 32'd1065666785;
      119: s256 = 32'd1067199482;
      120: s256 = 32'd1068571463;
      121: s256 = 32'd1069782521;
      122: s256 = 32'd1070832474;
      123: s256 = 32'd1071721163;
      124: s256 = 32'd1072448454;
      125: s256 = 32'd1073014239;
      126: s256 = 32'd1073418433;
      127: s256 = 32'd1073660973;
      128: s256 = 32'd1073741824;
      129: s256 = 32'd1073660973;
      130: s256 = 32'd1073418433;
      131: s256 = 32'd1073014239;
      132: s256 = 32'd1072448454;
      133: s256 = 32'd1071721163;
      134: s256 = 32'd1070832474;
      135: s256 = 32'd1069782521;
      136: s256 = 32'd1068571463;
      137: s256 = 32'd1067199482;
      138: s256 = 32'd1065666785;
      139: s256 = 32'd1063973603;
      140: s256 = 32'd1062120190;
      141: s256 = 32'd1060106825;
      142: s256 = 32'd1057933812;
      143: s256 = 32'd1055601479;
      144: s256 = 32'd1053110175;
      145: s256 = 32'd1050460278;
      146: s256 = 32'd1047652184;
      147: s256 = 32'd1044686318;
      148: s256 = 32'd1041563127;
      149: s256 = 32'd1038283079;
      150: s256 = 32'd1034846670;
      151: s256 = 32'd1031254417;
      152: s256 = 32'd1027506861;
      153: s256 = 32'd1023604566;
      154: s256 = 32'd1019548120;
      155: s256 = 32'd1015338134;
      156: s256 = 32'd1010975241;
      157: s256 = 32'd1006460100;
      158: s256 = 32'd1001793389;
      159: s256 = 32'd996975812;
      160: s256 = 32'd992008094;
      161: s256 = 32'd986890983;
      162: s256 = 32'd981625250;
      163: s256 = 32'd976211688;
      164: s256 = 32'd970651112;
      165: s256 = 32'd964944359;
      166: s256 = 32'd959092290;
      167: s256 = 32'd953095785;
      168: s256 = 32'd946955747;
      169: s256 = 32'd940673100;
      170: s256 = 32'd934248792;
      171: s256 = 32'd927683790;
      172: s256 = 32'd920979082;
      173: s256 = 32'd914135677;
      174: s256 = 32'd907154608;
      175: s256 = 32'd900036924;
      176: s256 = 32'd892783698;
      177: s256 = 32'd885396022;
      178: s256 = 32'd877875008;
      179: s256 = 32'd870221790;
      180: s256 = 32'd862437519;
      181: s256 = 32'd854523369;
      182: s256 = 32'd846480531;
      183: s256 = 32'd838310215;
      184: s256 = 32'd830013654;
      185: s256 = 32'd821592095;
      186: s256 = 32'd813046807;
      187: s256 = 32'd804379078;
      188: s256 = 32'd795590212;
      189: s256 = 32'd786681534;
      190: s256 = 32'd777654383;
      191: s256 = 32'd768510121;
      192: s256 = 32'd759250124;
      193: s256 = 32'd749875787;
      194: s256 = 32'd740388522;
      195: s256 = 32'd730789756;
      196: s256 = 32'd721080937;
      197: s256 = 32'd711263525;
      198: s256 = 32'd701338999;
      199: s256 = 32'd691308855;
      200: s256 = 32'd681174602;
      201: s256 = 32'd670937766;
      202: s256 = 32'd660599890;
      203: s256 = 32'd650162530;
      204: s256 = 32'd639627257;
      205: s256 = 32'd628995659;
      206: s256 = 32'd618269337;
      207: s256 = 32'd607449906;
      208: s256 = 32'd596538995;
      209: s256 = 32'd585538247;
      210: s256 = 32'd574449320;
      211: s256 = 32'd563273882;
      212: s256 = 32'd552013618;
      213: s256 = 32'd540670222;
      214: s256 = 32'd529245403;
      215: s256 = 32'd517740882;
      216: s256 = 32'd506158392;
      217: s256 = 32'd494499675;
      218: s256 = 32'd482766489;
      219: s256 = 32'd470960600;
      220: s256 = 32'd459083785;
      221: s256 = 32'd447137835;
      222: s256 = 32'd435124547;
      223: s256 = 32'd423045731;
      224: s256 = 32'd410903206;
      225: s256 = 32'd398698801;
      226: s256 = 32'd386434352;
      227: s256 = 32'd374111709;
      228: s256 = 32'd361732725;
      229: s256 = 32'd349299266;
      230: s256 = 32'd336813204;
      231: s256 = 32'd324276418;
      232: s256 = 32'd311690798;
      233: s256 = 32'd299058239;
      234: s256 = 32'd286380642;
      235: s256 = 32'd273659918;
      236: s256 = 32'd260897981;
      237: s256 = 32'd248096754;
      238: s256 = 32'd235258165;
      239: s256 = 32'd222384146;
      240: s256 = 32'd209476638;
      241: s256 = 32'd196537583;
      242: s256 = 32'd183568930;
      243: s256 = 32'd170572632;
      244: s256 = 32'd157550647;
      245: s256 = 32'd144504935;
      246: s256 = 32'd131437461;
      247: s256 = 32'd118350193;
      248: s256 = 32'd105245103;
      249: s256 = 32'd92124162;
      250: s256 = 32'd78989348;
      251: s256 = 32'd65842639;
      252: s256 = 32'd52686014;
      253: s256 = 32'd39521454;
      254: s256 = 32'd26350943;
      255: s256 = 32'd13176463;
    endcase
  always @(*)
    case(s526)
      0: s263 = 32'd1073741824;
      1: s263 = 32'd992008094;
      2: s263 = 32'd759250124;
      3: s263 = 32'd410903206;
      4: s263 = 32'd0;
      5: s263 = 32'd3884064090;
      6: s263 = 32'd3535717172;
      7: s263 = 32'd3302959202;
    endcase
  always @(*)
    case(s257)
      0: s277 = 32'd0;
      1: s277 = 32'd105245103;
      2: s277 = 32'd209476638;
      3: s277 = 32'd311690798;
      4: s277 = 32'd410903206;
      5: s277 = 32'd506158392;
      6: s277 = 32'd596538995;
      7: s277 = 32'd681174602;
      8: s277 = 32'd759250124;
      9: s277 = 32'd830013654;
      10: s277 = 32'd892783698;
      11: s277 = 32'd946955747;
      12: s277 = 32'd992008094;
      13: s277 = 32'd1027506861;
      14: s277 = 32'd1053110175;
      15: s277 = 32'd1068571463;
      16: s277 = 32'd1073741824;
      17: s277 = 32'd1068571463;
      18: s277 = 32'd1053110175;
      19: s277 = 32'd1027506861;
      20: s277 = 32'd992008094;
      21: s277 = 32'd946955747;
      22: s277 = 32'd892783698;
      23: s277 = 32'd830013654;
      24: s277 = 32'd759250124;
      25: s277 = 32'd681174602;
      26: s277 = 32'd596538995;
      27: s277 = 32'd506158392;
      28: s277 = 32'd410903206;
      29: s277 = 32'd311690798;
      30: s277 = 32'd209476638;
      31: s277 = 32'd105245103;
    endcase
  always @(*)
    case(s435)
      0: s525 = 32'd1073741824;
      1: s525 = 32'd1073721611;
      2: s525 = 32'd1073660973;
      3: s525 = 32'd1073559912;
      4: s525 = 32'd1073418433;
      5: s525 = 32'd1073236539;
      6: s525 = 32'd1073014239;
      7: s525 = 32'd1072751541;
      8: s525 = 32'd1072448454;
      9: s525 = 32'd1072104991;
      10: s525 = 32'd1071721163;
      11: s525 = 32'd1071296985;
      12: s525 = 32'd1070832474;
      13: s525 = 32'd1070327646;
      14: s525 = 32'd1069782521;
      15: s525 = 32'd1069197119;
      16: s525 = 32'd1068571463;
      17: s525 = 32'd1067905576;
      18: s525 = 32'd1067199482;
      19: s525 = 32'd1066453209;
      20: s525 = 32'd1065666785;
      21: s525 = 32'd1064840239;
      22: s525 = 32'd1063973603;
      23: s525 = 32'd1063066908;
      24: s525 = 32'd1062120190;
      25: s525 = 32'd1061133483;
      26: s525 = 32'd1060106825;
      27: s525 = 32'd1059040255;
      28: s525 = 32'd1057933812;
      29: s525 = 32'd1056787539;
      30: s525 = 32'd1055601479;
      31: s525 = 32'd1054375675;
      32: s525 = 32'd1053110175;
      33: s525 = 32'd1051805026;
      34: s525 = 32'd1050460278;
      35: s525 = 32'd1049075979;
      36: s525 = 32'd1047652184;
      37: s525 = 32'd1046188946;
      38: s525 = 32'd1044686318;
      39: s525 = 32'd1043144359;
      40: s525 = 32'd1041563127;
      41: s525 = 32'd1039942680;
      42: s525 = 32'd1038283079;
      43: s525 = 32'd1036584388;
      44: s525 = 32'd1034846670;
      45: s525 = 32'd1033069991;
      46: s525 = 32'd1031254417;
      47: s525 = 32'd1029400017;
      48: s525 = 32'd1027506861;
      49: s525 = 32'd1025575020;
      50: s525 = 32'd1023604566;
      51: s525 = 32'd1021595574;
      52: s525 = 32'd1019548120;
      53: s525 = 32'd1017462280;
      54: s525 = 32'd1015338134;
      55: s525 = 32'd1013175760;
      56: s525 = 32'd1010975241;
      57: s525 = 32'd1008736660;
      58: s525 = 32'd1006460100;
      59: s525 = 32'd1004145647;
      60: s525 = 32'd1001793389;
      61: s525 = 32'd999403414;
      62: s525 = 32'd996975812;
      63: s525 = 32'd994510674;
      64: s525 = 32'd992008094;
      65: s525 = 32'd989468165;
      66: s525 = 32'd986890983;
      67: s525 = 32'd984276645;
      68: s525 = 32'd981625250;
      69: s525 = 32'd978936897;
      70: s525 = 32'd976211688;
      71: s525 = 32'd973449725;
      72: s525 = 32'd970651112;
      73: s525 = 32'd967815955;
      74: s525 = 32'd964944359;
      75: s525 = 32'd962036435;
      76: s525 = 32'd959092290;
      77: s525 = 32'd956112036;
      78: s525 = 32'd953095785;
      79: s525 = 32'd950043650;
      80: s525 = 32'd946955747;
      81: s525 = 32'd943832191;
      82: s525 = 32'd940673100;
      83: s525 = 32'd937478594;
      84: s525 = 32'd934248792;
      85: s525 = 32'd930983817;
      86: s525 = 32'd927683790;
      87: s525 = 32'd924348836;
      88: s525 = 32'd920979082;
      89: s525 = 32'd917574653;
      90: s525 = 32'd914135677;
      91: s525 = 32'd910662286;
      92: s525 = 32'd907154608;
      93: s525 = 32'd903612776;
      94: s525 = 32'd900036924;
      95: s525 = 32'd896427186;
      96: s525 = 32'd892783698;
      97: s525 = 32'd889106597;
      98: s525 = 32'd885396022;
      99: s525 = 32'd881652112;
      100: s525 = 32'd877875008;
      101: s525 = 32'd874064853;
      102: s525 = 32'd870221790;
      103: s525 = 32'd866345963;
      104: s525 = 32'd862437519;
      105: s525 = 32'd858496605;
      106: s525 = 32'd854523369;
      107: s525 = 32'd850517961;
      108: s525 = 32'd846480531;
      109: s525 = 32'd842411231;
      110: s525 = 32'd838310215;
      111: s525 = 32'd834177638;
      112: s525 = 32'd830013654;
      113: s525 = 32'd825818420;
      114: s525 = 32'd821592095;
      115: s525 = 32'd817334837;
      116: s525 = 32'd813046807;
      117: s525 = 32'd808728167;
      118: s525 = 32'd804379078;
      119: s525 = 32'd799999705;
      120: s525 = 32'd795590212;
      121: s525 = 32'd791150766;
      122: s525 = 32'd786681534;
      123: s525 = 32'd782182683;
      124: s525 = 32'd777654383;
      125: s525 = 32'd773096806;
      126: s525 = 32'd768510121;
      127: s525 = 32'd763894503;
      128: s525 = 32'd759250124;
      129: s525 = 32'd754577161;
      130: s525 = 32'd749875787;
      131: s525 = 32'd745146182;
      132: s525 = 32'd740388522;
      133: s525 = 32'd735602987;
      134: s525 = 32'd730789756;
      135: s525 = 32'd725949012;
      136: s525 = 32'd721080937;
      137: s525 = 32'd716185713;
      138: s525 = 32'd711263525;
      139: s525 = 32'd706314558;
      140: s525 = 32'd701338999;
      141: s525 = 32'd696337035;
      142: s525 = 32'd691308855;
      143: s525 = 32'd686254647;
      144: s525 = 32'd681174602;
      145: s525 = 32'd676068911;
      146: s525 = 32'd670937766;
      147: s525 = 32'd665781361;
      148: s525 = 32'd660599890;
      149: s525 = 32'd655393547;
      150: s525 = 32'd650162530;
      151: s525 = 32'd644907034;
      152: s525 = 32'd639627257;
      153: s525 = 32'd634323399;
      154: s525 = 32'd628995659;
      155: s525 = 32'd623644238;
      156: s525 = 32'd618269337;
      157: s525 = 32'd612871159;
      158: s525 = 32'd607449906;
      159: s525 = 32'd602005783;
      160: s525 = 32'd596538995;
      161: s525 = 32'd591049747;
      162: s525 = 32'd585538247;
      163: s525 = 32'd580004702;
      164: s525 = 32'd574449320;
      165: s525 = 32'd568872310;
      166: s525 = 32'd563273882;
      167: s525 = 32'd557654248;
      168: s525 = 32'd552013618;
      169: s525 = 32'd546352205;
      170: s525 = 32'd540670222;
      171: s525 = 32'd534967883;
      172: s525 = 32'd529245403;
      173: s525 = 32'd523502998;
      174: s525 = 32'd517740882;
      175: s525 = 32'd511959274;
      176: s525 = 32'd506158392;
      177: s525 = 32'd500338452;
      178: s525 = 32'd494499675;
      179: s525 = 32'd488642280;
      180: s525 = 32'd482766489;
      181: s525 = 32'd476872521;
      182: s525 = 32'd470960600;
      183: s525 = 32'd465030947;
      184: s525 = 32'd459083785;
      185: s525 = 32'd453119340;
      186: s525 = 32'd447137835;
      187: s525 = 32'd441139495;
      188: s525 = 32'd435124547;
      189: s525 = 32'd429093217;
      190: s525 = 32'd423045731;
      191: s525 = 32'd416982318;
      192: s525 = 32'd410903206;
      193: s525 = 32'd404808624;
      194: s525 = 32'd398698801;
      195: s525 = 32'd392573967;
      196: s525 = 32'd386434352;
      197: s525 = 32'd380280189;
      198: s525 = 32'd374111709;
      199: s525 = 32'd367929143;
      200: s525 = 32'd361732725;
      201: s525 = 32'd355522688;
      202: s525 = 32'd349299266;
      203: s525 = 32'd343062693;
      204: s525 = 32'd336813204;
      205: s525 = 32'd330551034;
      206: s525 = 32'd324276418;
      207: s525 = 32'd317989594;
      208: s525 = 32'd311690798;
      209: s525 = 32'd305380267;
      210: s525 = 32'd299058239;
      211: s525 = 32'd292724951;
      212: s525 = 32'd286380642;
      213: s525 = 32'd280025551;
      214: s525 = 32'd273659918;
      215: s525 = 32'd267283981;
      216: s525 = 32'd260897981;
      217: s525 = 32'd254502159;
      218: s525 = 32'd248096754;
      219: s525 = 32'd241682009;
      220: s525 = 32'd235258165;
      221: s525 = 32'd228825463;
      222: s525 = 32'd222384146;
      223: s525 = 32'd215934457;
      224: s525 = 32'd209476638;
      225: s525 = 32'd203010932;
      226: s525 = 32'd196537583;
      227: s525 = 32'd190056834;
      228: s525 = 32'd183568930;
      229: s525 = 32'd177074114;
      230: s525 = 32'd170572632;
      231: s525 = 32'd164064728;
      232: s525 = 32'd157550647;
      233: s525 = 32'd151030634;
      234: s525 = 32'd144504935;
      235: s525 = 32'd137973795;
      236: s525 = 32'd131437461;
      237: s525 = 32'd124896178;
      238: s525 = 32'd118350193;
      239: s525 = 32'd111799753;
      240: s525 = 32'd105245103;
      241: s525 = 32'd98686490;
      242: s525 = 32'd92124162;
      243: s525 = 32'd85558366;
      244: s525 = 32'd78989348;
      245: s525 = 32'd72417357;
      246: s525 = 32'd65842639;
      247: s525 = 32'd59265442;
      248: s525 = 32'd52686014;
      249: s525 = 32'd46104602;
      250: s525 = 32'd39521454;
      251: s525 = 32'd32936819;
      252: s525 = 32'd26350943;
      253: s525 = 32'd19764075;
      254: s525 = 32'd13176463;
      255: s525 = 32'd6588355;
      256: s525 = 32'd0;
      257: s525 = 32'd4288378941;
      258: s525 = 32'd4281790833;
      259: s525 = 32'd4275203221;
      260: s525 = 32'd4268616353;
      261: s525 = 32'd4262030477;
      262: s525 = 32'd4255445842;
      263: s525 = 32'd4248862694;
      264: s525 = 32'd4242281282;
      265: s525 = 32'd4235701854;
      266: s525 = 32'd4229124657;
      267: s525 = 32'd4222549939;
      268: s525 = 32'd4215977948;
      269: s525 = 32'd4209408930;
      270: s525 = 32'd4202843134;
      271: s525 = 32'd4196280806;
      272: s525 = 32'd4189722193;
      273: s525 = 32'd4183167543;
      274: s525 = 32'd4176617103;
      275: s525 = 32'd4170071118;
      276: s525 = 32'd4163529835;
      277: s525 = 32'd4156993501;
      278: s525 = 32'd4150462361;
      279: s525 = 32'd4143936662;
      280: s525 = 32'd4137416649;
      281: s525 = 32'd4130902568;
      282: s525 = 32'd4124394664;
      283: s525 = 32'd4117893182;
      284: s525 = 32'd4111398366;
      285: s525 = 32'd4104910462;
      286: s525 = 32'd4098429713;
      287: s525 = 32'd4091956364;
      288: s525 = 32'd4085490658;
      289: s525 = 32'd4079032839;
      290: s525 = 32'd4072583150;
      291: s525 = 32'd4066141833;
      292: s525 = 32'd4059709131;
      293: s525 = 32'd4053285287;
      294: s525 = 32'd4046870542;
      295: s525 = 32'd4040465137;
      296: s525 = 32'd4034069315;
      297: s525 = 32'd4027683315;
      298: s525 = 32'd4021307378;
      299: s525 = 32'd4014941745;
      300: s525 = 32'd4008586654;
      301: s525 = 32'd4002242345;
      302: s525 = 32'd3995909057;
      303: s525 = 32'd3989587029;
      304: s525 = 32'd3983276498;
      305: s525 = 32'd3976977702;
      306: s525 = 32'd3970690878;
      307: s525 = 32'd3964416262;
      308: s525 = 32'd3958154092;
      309: s525 = 32'd3951904603;
      310: s525 = 32'd3945668030;
      311: s525 = 32'd3939444608;
      312: s525 = 32'd3933234571;
      313: s525 = 32'd3927038153;
      314: s525 = 32'd3920855587;
      315: s525 = 32'd3914687107;
      316: s525 = 32'd3908532944;
      317: s525 = 32'd3902393329;
      318: s525 = 32'd3896268495;
      319: s525 = 32'd3890158672;
      320: s525 = 32'd3884064090;
      321: s525 = 32'd3877984978;
      322: s525 = 32'd3871921565;
      323: s525 = 32'd3865874079;
      324: s525 = 32'd3859842749;
      325: s525 = 32'd3853827801;
      326: s525 = 32'd3847829461;
      327: s525 = 32'd3841847956;
      328: s525 = 32'd3835883511;
      329: s525 = 32'd3829936349;
      330: s525 = 32'd3824006696;
      331: s525 = 32'd3818094775;
      332: s525 = 32'd3812200807;
      333: s525 = 32'd3806325016;
      334: s525 = 32'd3800467621;
      335: s525 = 32'd3794628844;
      336: s525 = 32'd3788808904;
      337: s525 = 32'd3783008022;
      338: s525 = 32'd3777226414;
      339: s525 = 32'd3771464298;
      340: s525 = 32'd3765721893;
      341: s525 = 32'd3759999413;
      342: s525 = 32'd3754297074;
      343: s525 = 32'd3748615091;
      344: s525 = 32'd3742953678;
      345: s525 = 32'd3737313048;
      346: s525 = 32'd3731693414;
      347: s525 = 32'd3726094986;
      348: s525 = 32'd3720517976;
      349: s525 = 32'd3714962594;
      350: s525 = 32'd3709429049;
      351: s525 = 32'd3703917549;
      352: s525 = 32'd3698428301;
      353: s525 = 32'd3692961513;
      354: s525 = 32'd3687517390;
      355: s525 = 32'd3682096137;
      356: s525 = 32'd3676697959;
      357: s525 = 32'd3671323058;
      358: s525 = 32'd3665971637;
      359: s525 = 32'd3660643897;
      360: s525 = 32'd3655340039;
      361: s525 = 32'd3650060262;
      362: s525 = 32'd3644804766;
      363: s525 = 32'd3639573749;
      364: s525 = 32'd3634367406;
      365: s525 = 32'd3629185935;
      366: s525 = 32'd3624029530;
      367: s525 = 32'd3618898385;
      368: s525 = 32'd3613792694;
      369: s525 = 32'd3608712649;
      370: s525 = 32'd3603658441;
      371: s525 = 32'd3598630261;
      372: s525 = 32'd3593628297;
      373: s525 = 32'd3588652738;
      374: s525 = 32'd3583703771;
      375: s525 = 32'd3578781583;
      376: s525 = 32'd3573886359;
      377: s525 = 32'd3569018284;
      378: s525 = 32'd3564177540;
      379: s525 = 32'd3559364309;
      380: s525 = 32'd3554578774;
      381: s525 = 32'd3549821114;
      382: s525 = 32'd3545091509;
      383: s525 = 32'd3540390135;
      384: s525 = 32'd3535717172;
      385: s525 = 32'd3531072793;
      386: s525 = 32'd3526457175;
      387: s525 = 32'd3521870490;
      388: s525 = 32'd3517312913;
      389: s525 = 32'd3512784613;
      390: s525 = 32'd3508285762;
      391: s525 = 32'd3503816530;
      392: s525 = 32'd3499377084;
      393: s525 = 32'd3494967591;
      394: s525 = 32'd3490588218;
      395: s525 = 32'd3486239129;
      396: s525 = 32'd3481920489;
      397: s525 = 32'd3477632459;
      398: s525 = 32'd3473375201;
      399: s525 = 32'd3469148876;
      400: s525 = 32'd3464953642;
      401: s525 = 32'd3460789658;
      402: s525 = 32'd3456657081;
      403: s525 = 32'd3452556065;
      404: s525 = 32'd3448486765;
      405: s525 = 32'd3444449335;
      406: s525 = 32'd3440443927;
      407: s525 = 32'd3436470691;
      408: s525 = 32'd3432529777;
      409: s525 = 32'd3428621333;
      410: s525 = 32'd3424745506;
      411: s525 = 32'd3420902443;
      412: s525 = 32'd3417092288;
      413: s525 = 32'd3413315184;
      414: s525 = 32'd3409571274;
      415: s525 = 32'd3405860699;
      416: s525 = 32'd3402183598;
      417: s525 = 32'd3398540110;
      418: s525 = 32'd3394930372;
      419: s525 = 32'd3391354520;
      420: s525 = 32'd3387812688;
      421: s525 = 32'd3384305010;
      422: s525 = 32'd3380831619;
      423: s525 = 32'd3377392643;
      424: s525 = 32'd3373988214;
      425: s525 = 32'd3370618460;
      426: s525 = 32'd3367283506;
      427: s525 = 32'd3363983479;
      428: s525 = 32'd3360718504;
      429: s525 = 32'd3357488702;
      430: s525 = 32'd3354294196;
      431: s525 = 32'd3351135105;
      432: s525 = 32'd3348011549;
      433: s525 = 32'd3344923646;
      434: s525 = 32'd3341871511;
      435: s525 = 32'd3338855260;
      436: s525 = 32'd3335875006;
      437: s525 = 32'd3332930861;
      438: s525 = 32'd3330022937;
      439: s525 = 32'd3327151341;
      440: s525 = 32'd3324316184;
      441: s525 = 32'd3321517571;
      442: s525 = 32'd3318755608;
      443: s525 = 32'd3316030399;
      444: s525 = 32'd3313342046;
      445: s525 = 32'd3310690651;
      446: s525 = 32'd3308076313;
      447: s525 = 32'd3305499131;
      448: s525 = 32'd3302959202;
      449: s525 = 32'd3300456622;
      450: s525 = 32'd3297991484;
      451: s525 = 32'd3295563882;
      452: s525 = 32'd3293173907;
      453: s525 = 32'd3290821649;
      454: s525 = 32'd3288507196;
      455: s525 = 32'd3286230636;
      456: s525 = 32'd3283992055;
      457: s525 = 32'd3281791536;
      458: s525 = 32'd3279629162;
      459: s525 = 32'd3277505016;
      460: s525 = 32'd3275419176;
      461: s525 = 32'd3273371722;
      462: s525 = 32'd3271362730;
      463: s525 = 32'd3269392276;
      464: s525 = 32'd3267460435;
      465: s525 = 32'd3265567279;
      466: s525 = 32'd3263712879;
      467: s525 = 32'd3261897305;
      468: s525 = 32'd3260120626;
      469: s525 = 32'd3258382908;
      470: s525 = 32'd3256684217;
      471: s525 = 32'd3255024616;
      472: s525 = 32'd3253404169;
      473: s525 = 32'd3251822937;
      474: s525 = 32'd3250280978;
      475: s525 = 32'd3248778350;
      476: s525 = 32'd3247315112;
      477: s525 = 32'd3245891317;
      478: s525 = 32'd3244507018;
      479: s525 = 32'd3243162270;
      480: s525 = 32'd3241857121;
      481: s525 = 32'd3240591621;
      482: s525 = 32'd3239365817;
      483: s525 = 32'd3238179757;
      484: s525 = 32'd3237033484;
      485: s525 = 32'd3235927041;
      486: s525 = 32'd3234860471;
      487: s525 = 32'd3233833813;
      488: s525 = 32'd3232847106;
      489: s525 = 32'd3231900388;
      490: s525 = 32'd3230993693;
      491: s525 = 32'd3230127057;
      492: s525 = 32'd3229300511;
      493: s525 = 32'd3228514087;
      494: s525 = 32'd3227767814;
      495: s525 = 32'd3227061720;
      496: s525 = 32'd3226395833;
      497: s525 = 32'd3225770177;
      498: s525 = 32'd3225184775;
      499: s525 = 32'd3224639650;
      500: s525 = 32'd3224134822;
      501: s525 = 32'd3223670311;
      502: s525 = 32'd3223246133;
      503: s525 = 32'd3222862305;
      504: s525 = 32'd3222518842;
      505: s525 = 32'd3222215755;
      506: s525 = 32'd3221953057;
      507: s525 = 32'd3221730757;
      508: s525 = 32'd3221548863;
      509: s525 = 32'd3221407384;
      510: s525 = 32'd3221306323;
      511: s525 = 32'd3221245685;
    endcase
  always @(*)
    case(s681)
      0: s568 = 32'd1073741824;
      1: s568 = 32'd1072448454;
      2: s568 = 32'd1068571463;
      3: s568 = 32'd1062120190;
      4: s568 = 32'd1053110175;
      5: s568 = 32'd1041563127;
      6: s568 = 32'd1027506861;
      7: s568 = 32'd1010975241;
      8: s568 = 32'd992008094;
      9: s568 = 32'd970651112;
      10: s568 = 32'd946955747;
      11: s568 = 32'd920979082;
      12: s568 = 32'd892783698;
      13: s568 = 32'd862437519;
      14: s568 = 32'd830013654;
      15: s568 = 32'd795590212;
      16: s568 = 32'd759250124;
      17: s568 = 32'd721080937;
      18: s568 = 32'd681174602;
      19: s568 = 32'd639627257;
      20: s568 = 32'd596538995;
      21: s568 = 32'd552013618;
      22: s568 = 32'd506158392;
      23: s568 = 32'd459083785;
      24: s568 = 32'd410903206;
      25: s568 = 32'd361732725;
      26: s568 = 32'd311690798;
      27: s568 = 32'd260897981;
      28: s568 = 32'd209476638;
      29: s568 = 32'd157550647;
      30: s568 = 32'd105245103;
      31: s568 = 32'd52686014;
      32: s568 = 32'd0;
      33: s568 = 32'd4242281282;
      34: s568 = 32'd4189722193;
      35: s568 = 32'd4137416649;
      36: s568 = 32'd4085490658;
      37: s568 = 32'd4034069315;
      38: s568 = 32'd3983276498;
      39: s568 = 32'd3933234571;
      40: s568 = 32'd3884064090;
      41: s568 = 32'd3835883511;
      42: s568 = 32'd3788808904;
      43: s568 = 32'd3742953678;
      44: s568 = 32'd3698428301;
      45: s568 = 32'd3655340039;
      46: s568 = 32'd3613792694;
      47: s568 = 32'd3573886359;
      48: s568 = 32'd3535717172;
      49: s568 = 32'd3499377084;
      50: s568 = 32'd3464953642;
      51: s568 = 32'd3432529777;
      52: s568 = 32'd3402183598;
      53: s568 = 32'd3373988214;
      54: s568 = 32'd3348011549;
      55: s568 = 32'd3324316184;
      56: s568 = 32'd3302959202;
      57: s568 = 32'd3283992055;
      58: s568 = 32'd3267460435;
      59: s568 = 32'd3253404169;
      60: s568 = 32'd3241857121;
      61: s568 = 32'd3232847106;
      62: s568 = 32'd3226395833;
      63: s568 = 32'd3222518842;
    endcase
  always @(*)
    case(s305)
      0: s581 = 32'd0;
      1: s581 = 32'd26350943;
      2: s581 = 32'd52686014;
      3: s581 = 32'd78989348;
      4: s581 = 32'd105245103;
      5: s581 = 32'd131437461;
      6: s581 = 32'd157550647;
      7: s581 = 32'd183568930;
      8: s581 = 32'd209476638;
      9: s581 = 32'd235258165;
      10: s581 = 32'd260897981;
      11: s581 = 32'd286380642;
      12: s581 = 32'd311690798;
      13: s581 = 32'd336813204;
      14: s581 = 32'd361732725;
      15: s581 = 32'd386434352;
      16: s581 = 32'd410903206;
      17: s581 = 32'd435124547;
      18: s581 = 32'd459083785;
      19: s581 = 32'd482766489;
      20: s581 = 32'd506158392;
      21: s581 = 32'd529245403;
      22: s581 = 32'd552013618;
      23: s581 = 32'd574449320;
      24: s581 = 32'd596538995;
      25: s581 = 32'd618269337;
      26: s581 = 32'd639627257;
      27: s581 = 32'd660599890;
      28: s581 = 32'd681174602;
      29: s581 = 32'd701338999;
      30: s581 = 32'd721080937;
      31: s581 = 32'd740388522;
      32: s581 = 32'd759250124;
      33: s581 = 32'd777654383;
      34: s581 = 32'd795590212;
      35: s581 = 32'd813046807;
      36: s581 = 32'd830013654;
      37: s581 = 32'd846480531;
      38: s581 = 32'd862437519;
      39: s581 = 32'd877875008;
      40: s581 = 32'd892783698;
      41: s581 = 32'd907154608;
      42: s581 = 32'd920979082;
      43: s581 = 32'd934248792;
      44: s581 = 32'd946955747;
      45: s581 = 32'd959092290;
      46: s581 = 32'd970651112;
      47: s581 = 32'd981625250;
      48: s581 = 32'd992008094;
      49: s581 = 32'd1001793389;
      50: s581 = 32'd1010975241;
      51: s581 = 32'd1019548120;
      52: s581 = 32'd1027506861;
      53: s581 = 32'd1034846670;
      54: s581 = 32'd1041563127;
      55: s581 = 32'd1047652184;
      56: s581 = 32'd1053110175;
      57: s581 = 32'd1057933812;
      58: s581 = 32'd1062120190;
      59: s581 = 32'd1065666785;
      60: s581 = 32'd1068571463;
      61: s581 = 32'd1070832474;
      62: s581 = 32'd1072448454;
      63: s581 = 32'd1073418433;
      64: s581 = 32'd1073741824;
      65: s581 = 32'd1073418433;
      66: s581 = 32'd1072448454;
      67: s581 = 32'd1070832474;
      68: s581 = 32'd1068571463;
      69: s581 = 32'd1065666785;
      70: s581 = 32'd1062120190;
      71: s581 = 32'd1057933812;
      72: s581 = 32'd1053110175;
      73: s581 = 32'd1047652184;
      74: s581 = 32'd1041563127;
      75: s581 = 32'd1034846670;
      76: s581 = 32'd1027506861;
      77: s581 = 32'd1019548120;
      78: s581 = 32'd1010975241;
      79: s581 = 32'd1001793389;
      80: s581 = 32'd992008094;
      81: s581 = 32'd981625250;
      82: s581 = 32'd970651112;
      83: s581 = 32'd959092290;
      84: s581 = 32'd946955747;
      85: s581 = 32'd934248792;
      86: s581 = 32'd920979082;
      87: s581 = 32'd907154608;
      88: s581 = 32'd892783698;
      89: s581 = 32'd877875008;
      90: s581 = 32'd862437519;
      91: s581 = 32'd846480531;
      92: s581 = 32'd830013654;
      93: s581 = 32'd813046807;
      94: s581 = 32'd795590212;
      95: s581 = 32'd777654383;
      96: s581 = 32'd759250124;
      97: s581 = 32'd740388522;
      98: s581 = 32'd721080937;
      99: s581 = 32'd701338999;
      100: s581 = 32'd681174602;
      101: s581 = 32'd660599890;
      102: s581 = 32'd639627257;
      103: s581 = 32'd618269337;
      104: s581 = 32'd596538995;
      105: s581 = 32'd574449320;
      106: s581 = 32'd552013618;
      107: s581 = 32'd529245403;
      108: s581 = 32'd506158392;
      109: s581 = 32'd482766489;
      110: s581 = 32'd459083785;
      111: s581 = 32'd435124547;
      112: s581 = 32'd410903206;
      113: s581 = 32'd386434352;
      114: s581 = 32'd361732725;
      115: s581 = 32'd336813204;
      116: s581 = 32'd311690798;
      117: s581 = 32'd286380642;
      118: s581 = 32'd260897981;
      119: s581 = 32'd235258165;
      120: s581 = 32'd209476638;
      121: s581 = 32'd183568930;
      122: s581 = 32'd157550647;
      123: s581 = 32'd131437461;
      124: s581 = 32'd105245103;
      125: s581 = 32'd78989348;
      126: s581 = 32'd52686014;
      127: s581 = 32'd26350943;
    endcase
  always @(*)
    case(s310)
      0: s599 = s147;
      1: s599 = s138;
      2: s599 = s691;
      3: s599 = s20;
      4: s599 = s950;
      5: s599 = s864;
      6: s599 = s385;
      7: s599 = s271;
      default: s599 = s38;
    endcase
  always @(*)
    case(s406)
      0: s705 = s350;
      1: s705 = s674;
      2: s705 = 32'd0;
      3: s705 = s113;
    endcase
  always @(*)
    case(s406)
      0: s706 = s352;
      1: s706 = s676;
      2: s706 = 32'd0;
      3: s706 = s114;
    endcase
  always @(*)
    case(s305)
      0: s707 = 32'd1073741824;
      1: s707 = 32'd1073418433;
      2: s707 = 32'd1072448454;
      3: s707 = 32'd1070832474;
      4: s707 = 32'd1068571463;
      5: s707 = 32'd1065666785;
      6: s707 = 32'd1062120190;
      7: s707 = 32'd1057933812;
      8: s707 = 32'd1053110175;
      9: s707 = 32'd1047652184;
      10: s707 = 32'd1041563127;
      11: s707 = 32'd1034846670;
      12: s707 = 32'd1027506861;
      13: s707 = 32'd1019548120;
      14: s707 = 32'd1010975241;
      15: s707 = 32'd1001793389;
      16: s707 = 32'd992008094;
      17: s707 = 32'd981625250;
      18: s707 = 32'd970651112;
      19: s707 = 32'd959092290;
      20: s707 = 32'd946955747;
      21: s707 = 32'd934248792;
      22: s707 = 32'd920979082;
      23: s707 = 32'd907154608;
      24: s707 = 32'd892783698;
      25: s707 = 32'd877875008;
      26: s707 = 32'd862437519;
      27: s707 = 32'd846480531;
      28: s707 = 32'd830013654;
      29: s707 = 32'd813046807;
      30: s707 = 32'd795590212;
      31: s707 = 32'd777654383;
      32: s707 = 32'd759250124;
      33: s707 = 32'd740388522;
      34: s707 = 32'd721080937;
      35: s707 = 32'd701338999;
      36: s707 = 32'd681174602;
      37: s707 = 32'd660599890;
      38: s707 = 32'd639627257;
      39: s707 = 32'd618269337;
      40: s707 = 32'd596538995;
      41: s707 = 32'd574449320;
      42: s707 = 32'd552013618;
      43: s707 = 32'd529245403;
      44: s707 = 32'd506158392;
      45: s707 = 32'd482766489;
      46: s707 = 32'd459083785;
      47: s707 = 32'd435124547;
      48: s707 = 32'd410903206;
      49: s707 = 32'd386434352;
      50: s707 = 32'd361732725;
      51: s707 = 32'd336813204;
      52: s707 = 32'd311690798;
      53: s707 = 32'd286380642;
      54: s707 = 32'd260897981;
      55: s707 = 32'd235258165;
      56: s707 = 32'd209476638;
      57: s707 = 32'd183568930;
      58: s707 = 32'd157550647;
      59: s707 = 32'd131437461;
      60: s707 = 32'd105245103;
      61: s707 = 32'd78989348;
      62: s707 = 32'd52686014;
      63: s707 = 32'd26350943;
      64: s707 = 32'd0;
      65: s707 = 32'd4268616353;
      66: s707 = 32'd4242281282;
      67: s707 = 32'd4215977948;
      68: s707 = 32'd4189722193;
      69: s707 = 32'd4163529835;
      70: s707 = 32'd4137416649;
      71: s707 = 32'd4111398366;
      72: s707 = 32'd4085490658;
      73: s707 = 32'd4059709131;
      74: s707 = 32'd4034069315;
      75: s707 = 32'd4008586654;
      76: s707 = 32'd3983276498;
      77: s707 = 32'd3958154092;
      78: s707 = 32'd3933234571;
      79: s707 = 32'd3908532944;
      80: s707 = 32'd3884064090;
      81: s707 = 32'd3859842749;
      82: s707 = 32'd3835883511;
      83: s707 = 32'd3812200807;
      84: s707 = 32'd3788808904;
      85: s707 = 32'd3765721893;
      86: s707 = 32'd3742953678;
      87: s707 = 32'd3720517976;
      88: s707 = 32'd3698428301;
      89: s707 = 32'd3676697959;
      90: s707 = 32'd3655340039;
      91: s707 = 32'd3634367406;
      92: s707 = 32'd3613792694;
      93: s707 = 32'd3593628297;
      94: s707 = 32'd3573886359;
      95: s707 = 32'd3554578774;
      96: s707 = 32'd3535717172;
      97: s707 = 32'd3517312913;
      98: s707 = 32'd3499377084;
      99: s707 = 32'd3481920489;
      100: s707 = 32'd3464953642;
      101: s707 = 32'd3448486765;
      102: s707 = 32'd3432529777;
      103: s707 = 32'd3417092288;
      104: s707 = 32'd3402183598;
      105: s707 = 32'd3387812688;
      106: s707 = 32'd3373988214;
      107: s707 = 32'd3360718504;
      108: s707 = 32'd3348011549;
      109: s707 = 32'd3335875006;
      110: s707 = 32'd3324316184;
      111: s707 = 32'd3313342046;
      112: s707 = 32'd3302959202;
      113: s707 = 32'd3293173907;
      114: s707 = 32'd3283992055;
      115: s707 = 32'd3275419176;
      116: s707 = 32'd3267460435;
      117: s707 = 32'd3260120626;
      118: s707 = 32'd3253404169;
      119: s707 = 32'd3247315112;
      120: s707 = 32'd3241857121;
      121: s707 = 32'd3237033484;
      122: s707 = 32'd3232847106;
      123: s707 = 32'd3229300511;
      124: s707 = 32'd3226395833;
      125: s707 = 32'd3224134822;
      126: s707 = 32'd3222518842;
      127: s707 = 32'd3221548863;
    endcase
  always @(*)
    case(s76)
      0: s747 = 32'd1073741824;
      1: s747 = 32'd1073660973;
      2: s747 = 32'd1073418433;
      3: s747 = 32'd1073014239;
      4: s747 = 32'd1072448454;
      5: s747 = 32'd1071721163;
      6: s747 = 32'd1070832474;
      7: s747 = 32'd1069782521;
      8: s747 = 32'd1068571463;
      9: s747 = 32'd1067199482;
      10: s747 = 32'd1065666785;
      11: s747 = 32'd1063973603;
      12: s747 = 32'd1062120190;
      13: s747 = 32'd1060106825;
      14: s747 = 32'd1057933812;
      15: s747 = 32'd1055601479;
      16: s747 = 32'd1053110175;
      17: s747 = 32'd1050460278;
      18: s747 = 32'd1047652184;
      19: s747 = 32'd1044686318;
      20: s747 = 32'd1041563127;
      21: s747 = 32'd1038283079;
      22: s747 = 32'd1034846670;
      23: s747 = 32'd1031254417;
      24: s747 = 32'd1027506861;
      25: s747 = 32'd1023604566;
      26: s747 = 32'd1019548120;
      27: s747 = 32'd1015338134;
      28: s747 = 32'd1010975241;
      29: s747 = 32'd1006460100;
      30: s747 = 32'd1001793389;
      31: s747 = 32'd996975812;
      32: s747 = 32'd992008094;
      33: s747 = 32'd986890983;
      34: s747 = 32'd981625250;
      35: s747 = 32'd976211688;
      36: s747 = 32'd970651112;
      37: s747 = 32'd964944359;
      38: s747 = 32'd959092290;
      39: s747 = 32'd953095785;
      40: s747 = 32'd946955747;
      41: s747 = 32'd940673100;
      42: s747 = 32'd934248792;
      43: s747 = 32'd927683790;
      44: s747 = 32'd920979082;
      45: s747 = 32'd914135677;
      46: s747 = 32'd907154608;
      47: s747 = 32'd900036924;
      48: s747 = 32'd892783698;
      49: s747 = 32'd885396022;
      50: s747 = 32'd877875008;
      51: s747 = 32'd870221790;
      52: s747 = 32'd862437519;
      53: s747 = 32'd854523369;
      54: s747 = 32'd846480531;
      55: s747 = 32'd838310215;
      56: s747 = 32'd830013654;
      57: s747 = 32'd821592095;
      58: s747 = 32'd813046807;
      59: s747 = 32'd804379078;
      60: s747 = 32'd795590212;
      61: s747 = 32'd786681534;
      62: s747 = 32'd777654383;
      63: s747 = 32'd768510121;
      64: s747 = 32'd759250124;
      65: s747 = 32'd749875787;
      66: s747 = 32'd740388522;
      67: s747 = 32'd730789756;
      68: s747 = 32'd721080937;
      69: s747 = 32'd711263525;
      70: s747 = 32'd701338999;
      71: s747 = 32'd691308855;
      72: s747 = 32'd681174602;
      73: s747 = 32'd670937766;
      74: s747 = 32'd660599890;
      75: s747 = 32'd650162530;
      76: s747 = 32'd639627257;
      77: s747 = 32'd628995659;
      78: s747 = 32'd618269337;
      79: s747 = 32'd607449906;
      80: s747 = 32'd596538995;
      81: s747 = 32'd585538247;
      82: s747 = 32'd574449320;
      83: s747 = 32'd563273882;
      84: s747 = 32'd552013618;
      85: s747 = 32'd540670222;
      86: s747 = 32'd529245403;
      87: s747 = 32'd517740882;
      88: s747 = 32'd506158392;
      89: s747 = 32'd494499675;
      90: s747 = 32'd482766489;
      91: s747 = 32'd470960600;
      92: s747 = 32'd459083785;
      93: s747 = 32'd447137835;
      94: s747 = 32'd435124547;
      95: s747 = 32'd423045731;
      96: s747 = 32'd410903206;
      97: s747 = 32'd398698801;
      98: s747 = 32'd386434352;
      99: s747 = 32'd374111709;
      100: s747 = 32'd361732725;
      101: s747 = 32'd349299266;
      102: s747 = 32'd336813204;
      103: s747 = 32'd324276418;
      104: s747 = 32'd311690798;
      105: s747 = 32'd299058239;
      106: s747 = 32'd286380642;
      107: s747 = 32'd273659918;
      108: s747 = 32'd260897981;
      109: s747 = 32'd248096754;
      110: s747 = 32'd235258165;
      111: s747 = 32'd222384146;
      112: s747 = 32'd209476638;
      113: s747 = 32'd196537583;
      114: s747 = 32'd183568930;
      115: s747 = 32'd170572632;
      116: s747 = 32'd157550647;
      117: s747 = 32'd144504935;
      118: s747 = 32'd131437461;
      119: s747 = 32'd118350193;
      120: s747 = 32'd105245103;
      121: s747 = 32'd92124162;
      122: s747 = 32'd78989348;
      123: s747 = 32'd65842639;
      124: s747 = 32'd52686014;
      125: s747 = 32'd39521454;
      126: s747 = 32'd26350943;
      127: s747 = 32'd13176463;
      128: s747 = 32'd0;
      129: s747 = 32'd4281790833;
      130: s747 = 32'd4268616353;
      131: s747 = 32'd4255445842;
      132: s747 = 32'd4242281282;
      133: s747 = 32'd4229124657;
      134: s747 = 32'd4215977948;
      135: s747 = 32'd4202843134;
      136: s747 = 32'd4189722193;
      137: s747 = 32'd4176617103;
      138: s747 = 32'd4163529835;
      139: s747 = 32'd4150462361;
      140: s747 = 32'd4137416649;
      141: s747 = 32'd4124394664;
      142: s747 = 32'd4111398366;
      143: s747 = 32'd4098429713;
      144: s747 = 32'd4085490658;
      145: s747 = 32'd4072583150;
      146: s747 = 32'd4059709131;
      147: s747 = 32'd4046870542;
      148: s747 = 32'd4034069315;
      149: s747 = 32'd4021307378;
      150: s747 = 32'd4008586654;
      151: s747 = 32'd3995909057;
      152: s747 = 32'd3983276498;
      153: s747 = 32'd3970690878;
      154: s747 = 32'd3958154092;
      155: s747 = 32'd3945668030;
      156: s747 = 32'd3933234571;
      157: s747 = 32'd3920855587;
      158: s747 = 32'd3908532944;
      159: s747 = 32'd3896268495;
      160: s747 = 32'd3884064090;
      161: s747 = 32'd3871921565;
      162: s747 = 32'd3859842749;
      163: s747 = 32'd3847829461;
      164: s747 = 32'd3835883511;
      165: s747 = 32'd3824006696;
      166: s747 = 32'd3812200807;
      167: s747 = 32'd3800467621;
      168: s747 = 32'd3788808904;
      169: s747 = 32'd3777226414;
      170: s747 = 32'd3765721893;
      171: s747 = 32'd3754297074;
      172: s747 = 32'd3742953678;
      173: s747 = 32'd3731693414;
      174: s747 = 32'd3720517976;
      175: s747 = 32'd3709429049;
      176: s747 = 32'd3698428301;
      177: s747 = 32'd3687517390;
      178: s747 = 32'd3676697959;
      179: s747 = 32'd3665971637;
      180: s747 = 32'd3655340039;
      181: s747 = 32'd3644804766;
      182: s747 = 32'd3634367406;
      183: s747 = 32'd3624029530;
      184: s747 = 32'd3613792694;
      185: s747 = 32'd3603658441;
      186: s747 = 32'd3593628297;
      187: s747 = 32'd3583703771;
      188: s747 = 32'd3573886359;
      189: s747 = 32'd3564177540;
      190: s747 = 32'd3554578774;
      191: s747 = 32'd3545091509;
      192: s747 = 32'd3535717172;
      193: s747 = 32'd3526457175;
      194: s747 = 32'd3517312913;
      195: s747 = 32'd3508285762;
      196: s747 = 32'd3499377084;
      197: s747 = 32'd3490588218;
      198: s747 = 32'd3481920489;
      199: s747 = 32'd3473375201;
      200: s747 = 32'd3464953642;
      201: s747 = 32'd3456657081;
      202: s747 = 32'd3448486765;
      203: s747 = 32'd3440443927;
      204: s747 = 32'd3432529777;
      205: s747 = 32'd3424745506;
      206: s747 = 32'd3417092288;
      207: s747 = 32'd3409571274;
      208: s747 = 32'd3402183598;
      209: s747 = 32'd3394930372;
      210: s747 = 32'd3387812688;
      211: s747 = 32'd3380831619;
      212: s747 = 32'd3373988214;
      213: s747 = 32'd3367283506;
      214: s747 = 32'd3360718504;
      215: s747 = 32'd3354294196;
      216: s747 = 32'd3348011549;
      217: s747 = 32'd3341871511;
      218: s747 = 32'd3335875006;
      219: s747 = 32'd3330022937;
      220: s747 = 32'd3324316184;
      221: s747 = 32'd3318755608;
      222: s747 = 32'd3313342046;
      223: s747 = 32'd3308076313;
      224: s747 = 32'd3302959202;
      225: s747 = 32'd3297991484;
      226: s747 = 32'd3293173907;
      227: s747 = 32'd3288507196;
      228: s747 = 32'd3283992055;
      229: s747 = 32'd3279629162;
      230: s747 = 32'd3275419176;
      231: s747 = 32'd3271362730;
      232: s747 = 32'd3267460435;
      233: s747 = 32'd3263712879;
      234: s747 = 32'd3260120626;
      235: s747 = 32'd3256684217;
      236: s747 = 32'd3253404169;
      237: s747 = 32'd3250280978;
      238: s747 = 32'd3247315112;
      239: s747 = 32'd3244507018;
      240: s747 = 32'd3241857121;
      241: s747 = 32'd3239365817;
      242: s747 = 32'd3237033484;
      243: s747 = 32'd3234860471;
      244: s747 = 32'd3232847106;
      245: s747 = 32'd3230993693;
      246: s747 = 32'd3229300511;
      247: s747 = 32'd3227767814;
      248: s747 = 32'd3226395833;
      249: s747 = 32'd3225184775;
      250: s747 = 32'd3224134822;
      251: s747 = 32'd3223246133;
      252: s747 = 32'd3222518842;
      253: s747 = 32'd3221953057;
      254: s747 = 32'd3221548863;
      255: s747 = 32'd3221306323;
    endcase
  always @(*)
    case(s71)
      0: s797 = 32'd1073741824;
      1: s797 = 32'd1053110175;
      2: s797 = 32'd992008094;
      3: s797 = 32'd892783698;
      4: s797 = 32'd759250124;
      5: s797 = 32'd596538995;
      6: s797 = 32'd410903206;
      7: s797 = 32'd209476638;
      8: s797 = 32'd0;
      9: s797 = 32'd4085490658;
      10: s797 = 32'd3884064090;
      11: s797 = 32'd3698428301;
      12: s797 = 32'd3535717172;
      13: s797 = 32'd3402183598;
      14: s797 = 32'd3302959202;
      15: s797 = 32'd3241857121;
    endcase
  always @(*)
    case(s257)
      0: s804 = 32'd1073741824;
      1: s804 = 32'd1068571463;
      2: s804 = 32'd1053110175;
      3: s804 = 32'd1027506861;
      4: s804 = 32'd992008094;
      5: s804 = 32'd946955747;
      6: s804 = 32'd892783698;
      7: s804 = 32'd830013654;
      8: s804 = 32'd759250124;
      9: s804 = 32'd681174602;
      10: s804 = 32'd596538995;
      11: s804 = 32'd506158392;
      12: s804 = 32'd410903206;
      13: s804 = 32'd311690798;
      14: s804 = 32'd209476638;
      15: s804 = 32'd105245103;
      16: s804 = 32'd0;
      17: s804 = 32'd4189722193;
      18: s804 = 32'd4085490658;
      19: s804 = 32'd3983276498;
      20: s804 = 32'd3884064090;
      21: s804 = 32'd3788808904;
      22: s804 = 32'd3698428301;
      23: s804 = 32'd3613792694;
      24: s804 = 32'd3535717172;
      25: s804 = 32'd3464953642;
      26: s804 = 32'd3402183598;
      27: s804 = 32'd3348011549;
      28: s804 = 32'd3302959202;
      29: s804 = 32'd3267460435;
      30: s804 = 32'd3241857121;
      31: s804 = 32'd3226395833;
    endcase
  always @(*)
    case(s71)
      0: s809 = 32'd0;
      1: s809 = 32'd209476638;
      2: s809 = 32'd410903206;
      3: s809 = 32'd596538995;
      4: s809 = 32'd759250124;
      5: s809 = 32'd892783698;
      6: s809 = 32'd992008094;
      7: s809 = 32'd1053110175;
      8: s809 = 32'd1073741824;
      9: s809 = 32'd1053110175;
      10: s809 = 32'd992008094;
      11: s809 = 32'd892783698;
      12: s809 = 32'd759250124;
      13: s809 = 32'd596538995;
      14: s809 = 32'd410903206;
      15: s809 = 32'd209476638;
    endcase
  always @(*)
    case(s406)
      0: s890 = 32'd0;
      1: s890 = s676;
      2: s890 = s352;
      3: s890 = s676;
    endcase
  always @(*)
    case(s406)
      0: s891 = 32'd0;
      1: s891 = s674;
      2: s891 = s350;
      3: s891 = s674;
    endcase
  always @(*)
    case(s55)
      0: s944 = 9'd0;
      1: s944 = 9'd1;
      2: s944 = 9'd3;
      3: s944 = 9'd7;
      4: s944 = 9'd15;
      5: s944 = 9'd31;
      6: s944 = 9'd63;
      7: s944 = 9'd127;
      8: s944 = 9'd255;
      9: s944 = 9'd511;
      10: s944 = 9'd510;
      11: s944 = 9'd508;
      12: s944 = 9'd504;
      13: s944 = 9'd496;
      14: s944 = 9'd480;
      15: s944 = 9'd448;
      16: s944 = 9'd384;
      default: s944 = 9'd256;
    endcase
  always @(*)
    case(s681)
      0: s945 = 32'd0;
      1: s945 = 32'd52686014;
      2: s945 = 32'd105245103;
      3: s945 = 32'd157550647;
      4: s945 = 32'd209476638;
      5: s945 = 32'd260897981;
      6: s945 = 32'd311690798;
      7: s945 = 32'd361732725;
      8: s945 = 32'd410903206;
      9: s945 = 32'd459083785;
      10: s945 = 32'd506158392;
      11: s945 = 32'd552013618;
      12: s945 = 32'd596538995;
      13: s945 = 32'd639627257;
      14: s945 = 32'd681174602;
      15: s945 = 32'd721080937;
      16: s945 = 32'd759250124;
      17: s945 = 32'd795590212;
      18: s945 = 32'd830013654;
      19: s945 = 32'd862437519;
      20: s945 = 32'd892783698;
      21: s945 = 32'd920979082;
      22: s945 = 32'd946955747;
      23: s945 = 32'd970651112;
      24: s945 = 32'd992008094;
      25: s945 = 32'd1010975241;
      26: s945 = 32'd1027506861;
      27: s945 = 32'd1041563127;
      28: s945 = 32'd1053110175;
      29: s945 = 32'd1062120190;
      30: s945 = 32'd1068571463;
      31: s945 = 32'd1072448454;
      32: s945 = 32'd1073741824;
      33: s945 = 32'd1072448454;
      34: s945 = 32'd1068571463;
      35: s945 = 32'd1062120190;
      36: s945 = 32'd1053110175;
      37: s945 = 32'd1041563127;
      38: s945 = 32'd1027506861;
      39: s945 = 32'd1010975241;
      40: s945 = 32'd992008094;
      41: s945 = 32'd970651112;
      42: s945 = 32'd946955747;
      43: s945 = 32'd920979082;
      44: s945 = 32'd892783698;
      45: s945 = 32'd862437519;
      46: s945 = 32'd830013654;
      47: s945 = 32'd795590212;
      48: s945 = 32'd759250124;
      49: s945 = 32'd721080937;
      50: s945 = 32'd681174602;
      51: s945 = 32'd639627257;
      52: s945 = 32'd596538995;
      53: s945 = 32'd552013618;
      54: s945 = 32'd506158392;
      55: s945 = 32'd459083785;
      56: s945 = 32'd410903206;
      57: s945 = 32'd361732725;
      58: s945 = 32'd311690798;
      59: s945 = 32'd260897981;
      60: s945 = 32'd209476638;
      61: s945 = 32'd157550647;
      62: s945 = 32'd105245103;
      63: s945 = 32'd52686014;
    endcase
  always @(posedge clk)
    begin
      s4 [0] <= s543;
      for (i = 1; i < 20; i = i + 1)
        s4 [i] <= s4 [i - 1];
      s8 [s74] <= s570;
      s7 <= s8 [s369];
      s9 <= s24;
      s10 <= s234;
      s11 <= s395;
      s13 [0] <= s928;
      for (i = 1; i < 15; i = i + 1)
        s13 [i] <= s13 [i - 1];
      s14 <= s716;
      s15 <= s717;
      s17 [s762] <= s333;
      s16 <= s17 [s715];
      s18 <= s705;
      s19 <= s706;
      s23 [0] <= s344;
      for (i = 1; i < 30; i = i + 1)
        s23 [i] <= s23 [i - 1];
      s25 [s906] <= s833;
      s24 <= s25 [s418];
      s26 <= s290;
      s27 <= s649;
      s40 [0] <= s360;
      for (i = 1; i < 595; i = i + 1)
        s40 [i] <= s40 [i - 1];
      s41 <= s354;
      s42 <= s355;
      s45 <= s6;
      s46 <= s95;
      s47 <= s96;
      s49 [0] <= s252;
      for (i = 1; i < 137; i = i + 1)
        s49 [i] <= s49 [i - 1];
      s52 <= s447;
      s54 [s348] <= s941;
      s53 <= s54 [s510];
      s55 <= s316;
      s57 [0] <= s600;
      for (i = 1; i < 4; i = i + 1)
        s57 [i] <= s57 [i - 1];
      s59 [0] <= s601;
      for (i = 1; i < 4; i = i + 1)
        s59 [i] <= s59 [i - 1];
      s61 <= s934;
      s62 <= s935;
      s66 <= s295;
      s67 <= s296;
      s69 <= s809;
      s72 [0] <= s762;
      for (i = 1; i < 11; i = i + 1)
        s72 [i] <= s72 [i - 1];
      s75 [0] <= s369;
      for (i = 1; i < 7; i = i + 1)
        s75 [i] <= s75 [i - 1];
      s77 [0] <= s236;
      for (i = 1; i < 131; i = i + 1)
        s77 [i] <= s77 [i - 1];
      s78 <= s313;
      s82 <= s373;
      s84 [0] <= s865;
      for (i = 1; i < 4; i = i + 1)
        s84 [i] <= s84 [i - 1];
      s89 [0] <= s870;
      for (i = 1; i < 4; i = i + 1)
        s89 [i] <= s89 [i - 1];
      s90 <= s532;
      s92 [0] <= s748;
      for (i = 1; i < 4; i = i + 1)
        s92 [i] <= s92 [i - 1];
      s94 [0] <= s749;
      for (i = 1; i < 4; i = i + 1)
        s94 [i] <= s94 [i - 1];
      s104 <= s277;
      s106 <= s157;
      s107 <= s85;
      s110 <= s707;
      s113 <= s647;
      s114 <= s648;
      s116 [0] <= s168;
      for (i = 1; i < 3; i = i + 1)
        s116 [i] <= s116 [i - 1];
      s118 [0] <= s169;
      for (i = 1; i < 3; i = i + 1)
        s118 [i] <= s118 [i - 1];
      s119 <= s755;
      s120 <= s281;
      s126 [0] <= s370;
      for (i = 1; i < 3; i = i + 1)
        s126 [i] <= s126 [i - 1];
      s128 [0] <= s371;
      for (i = 1; i < 3; i = i + 1)
        s128 [i] <= s128 [i - 1];
      s129 <= s888;
      s130 <= s791;
      s132 <= s604;
      s133 <= s605;
      s135 [0] <= s735;
      for (i = 1; i < 3; i = i + 1)
        s135 [i] <= s135 [i - 1];
      s137 [0] <= s736;
      for (i = 1; i < 3; i = i + 1)
        s137 [i] <= s137 [i - 1];
      s140 <= s494;
      s143 <= s177;
      s144 <= s178;
      s146 <= s151;
      s148 [0] <= s348;
      for (i = 1; i < 9; i = i + 1)
        s148 [i] <= s148 [i - 1];
      s154 <= s539;
      s156 [0] <= s340;
      for (i = 1; i < 73; i = i + 1)
        s156 [i] <= s156 [i - 1];
      s158 [s460] <= s639;
      s157 <= s158 [s154];
      s161 <= s815;
      s162 <= s816;
      s164 <= s567;
      s165 <= s562;
      s175 <= s638;
      s176 <= s813;
      s180 <= s484;
      s181 <= s485;
      s186 <= s440;
      s189 <= s804;
      s190 <= s599;
      s192 [0] <= s257;
      for (i = 1; i < 270; i = i + 1)
        s192 [i] <= s192 [i - 1];
      s194 <= s53;
      s196 [s272] <= s585;
      s195 <= s196 [s255];
      s204 [s922] <= s911;
      s203 <= s204 [s524];
      s205 <= s314;
      s207 [0] <= s155;
      for (i = 1; i < 68; i = i + 1)
        s207 [i] <= s207 [i - 1];
      s208 <= s551;
      s209 <= s342;
      s210 <= s343;
      s213 [0] <= s30;
      for (i = 1; i < 4; i = i + 1)
        s213 [i] <= s213 [i - 1];
      s215 [0] <= s31;
      for (i = 1; i < 4; i = i + 1)
        s215 [i] <= s215 [i - 1];
      s220 <= s338;
      s222 [0] <= s239;
      for (i = 1; i < 255; i = i + 1)
        s222 [i] <= s222 [i - 1];
      s223 <= s87;
      s226 [0] <= s688;
      for (i = 1; i < 3; i = i + 1)
        s226 [i] <= s226 [i - 1];
      s228 [0] <= s689;
      for (i = 1; i < 3; i = i + 1)
        s228 [i] <= s228 [i - 1];
      s231 <= s806;
      s232 <= s840;
      s235 <= s859;
      s237 [0] <= s606;
      for (i = 1; i < 127; i = i + 1)
        s237 [i] <= s237 [i - 1];
      s239 <= s388;
      s241 [0] <= s392;
      for (i = 1; i < 6; i = i + 1)
        s241 [i] <= s241 [i - 1];
      s242 <= s919;
      s245 <= s592;
      s247 [0] <= s71;
      for (i = 1; i < 296; i = i + 1)
        s247 [i] <= s247 [i - 1];
      s251 [0] <= s356;
      for (i = 1; i < 15; i = i + 1)
        s251 [i] <= s251 [i - 1];
      s253 [0] <= s473;
      for (i = 1; i < 576; i = i + 1)
        s253 [i] <= s253 [i - 1];
      s254 <= s438;
      s255 <= s190;
      s258 [0] <= s508;
      for (i = 1; i < 19; i = i + 1)
        s258 [i] <= s258 [i - 1];
      s261 <= s920;
      s262 <= s921;
      s268 [s250] <= s708;
      s267 <= s268 [s356];
      s269 <= s443;
      s273 [0] <= s255;
      for (i = 1; i < 255; i = i + 1)
        s273 [i] <= s273 [i - 1];
      s274 <= s401;
      s275 <= s402;
      s276 <= s139;
      s278 <= s183;
      s280 [0] <= s530;
      for (i = 1; i < 30; i = i + 1)
        s280 [i] <= s280 [i - 1];
      s286 <= s364;
      s287 <= s365;
      s288 <= s760;
      s292 [0] <= s320;
      for (i = 1; i < 262; i = i + 1)
        s292 [i] <= s292 [i - 1];
      s294 <= s714;
      s297 <= s289;
      s300 [s718] <= s60;
      s299 <= s300 [s254];
      s302 [0] <= s386;
      for (i = 1; i < 4; i = i + 1)
        s302 [i] <= s302 [i - 1];
      s304 [0] <= s387;
      for (i = 1; i < 4; i = i + 1)
        s304 [i] <= s304 [i - 1];
      s306 [0] <= s737;
      for (i = 1; i < 67; i = i + 1)
        s306 [i] <= s306 [i - 1];
      s309 <= s552;
      s308 <= s309;
      s310 <= s283;
      s312 <= s331;
      s315 [s367] <= s167;
      s314 <= s315 [s832];
      s319 [0] <= s594;
      for (i = 1; i < 10; i = i + 1)
        s319 [i] <= s319 [i - 1];
      s321 [0] <= s802;
      for (i = 1; i < 4; i = i + 1)
        s321 [i] <= s321 [i - 1];
      s326 <= s449;
      s332 [s508] <= s166;
      s331 <= s332 [s884];
      s335 <= s468;
      s336 <= s939;
      s337 <= s216;
      s341 [0] <= s474;
      for (i = 1; i < 566; i = i + 1)
        s341 [i] <= s341 [i - 1];
      s347 [0] <= s458;
      for (i = 1; i < 10; i = i + 1)
        s347 [i] <= s347 [i - 1];
      s349 [0] <= s510;
      for (i = 1; i < 255; i = i + 1)
        s349 [i] <= s349 [i - 1];
      s351 [0] <= s698;
      for (i = 1; i < 3; i = i + 1)
        s351 [i] <= s351 [i - 1];
      s353 [0] <= s699;
      for (i = 1; i < 3; i = i + 1)
        s353 [i] <= s353 [i - 1];
      s356 <= s112;
      s357 <= s256;
      s361 <= s778;
      s366 <= s121;
      s368 [0] <= s832;
      for (i = 1; i < 31; i = i + 1)
        s368 [i] <= s368 [i - 1];
      s369 <= s105;
      s372 <= s326;
      s374 <= s598;
      s375 <= s383;
      s376 <= s152;
      s378 [0] <= s159;
      for (i = 1; i < 3; i = i + 1)
        s378 [i] <= s378 [i - 1];
      s380 [0] <= s160;
      for (i = 1; i < 3; i = i + 1)
        s380 [i] <= s380 [i - 1];
      s382 [0] <= s471;
      for (i = 1; i < 586; i = i + 1)
        s382 [i] <= s382 [i - 1];
      s384 <= s244;
      s389 <= s233;
      s390 <= s890;
      s391 <= s891;
      s393 [0] <= s702;
      for (i = 1; i < 6; i = i + 1)
        s393 [i] <= s393 [i - 1];
      s394 <= s767;
      s396 <= s779;
      s399 <= s577;
      s400 <= s578;
      s404 [0] <= s946;
      for (i = 1; i < 256; i = i + 1)
        s404 [i] <= s404 [i - 1];
      s405 <= s182;
      s407 [0] <= s288;
      for (i = 1; i < 10; i = i + 1)
        s407 [i] <= s407 [i - 1];
      s408 <= s267;
      s410 [s751] <= s709;
      s409 <= s410 [s107];
      s412 <= s285;
      s414 [0] <= s630;
      for (i = 1; i < 4; i = i + 1)
        s414 [i] <= s414 [i - 1];
      s416 [0] <= s631;
      for (i = 1; i < 4; i = i + 1)
        s416 [i] <= s416 [i - 1];
      s417 <= s86;
      s418 <= s431;
      s419 <= s428;
      s420 <= s634;
      s421 <= s179;
      s424 <= s21;
      s427 <= s810;
      s429 <= s264;
      s433 [s565] <= s122;
      s432 <= s433 [s417];
      s434 <= s263;
      s436 [0] <= s147;
      for (i = 1; i < 250; i = i + 1)
        s436 [i] <= s436 [i - 1];
      s439 <= s284;
      s440 <= s188;
      s442 [0] <= s528;
      for (i = 1; i < 4; i = i + 1)
        s442 [i] <= s442 [i - 1];
      s443 <= s163;
      s444 <= s448;
      s445 <= s73;
      s446 <= s282;
      s452 <= s729;
      s455 <= s298;
      s456 <= s949;
      s459 [0] <= s936;
      for (i = 1; i < 10; i = i + 1)
        s459 [i] <= s459 [i - 1];
      s461 [0] <= s154;
      for (i = 1; i < 3; i = i + 1)
        s461 [i] <= s461 [i - 1];
      s462 <= s195;
      s465 <= s79;
      s469 <= s563;
      s470 <= s564;
      s481 [0] <= s792;
      for (i = 1; i < 6; i = i + 1)
        s481 [i] <= s481 [i - 1];
      s483 [0] <= s793;
      for (i = 1; i < 6; i = i + 1)
        s483 [i] <= s483 [i - 1];
      s487 [0] <= s908;
      for (i = 1; i < 4; i = i + 1)
        s487 [i] <= s487 [i - 1];
      s489 [0] <= s909;
      for (i = 1; i < 4; i = i + 1)
        s489 [i] <= s489 [i - 1];
      s491 [0] <= s794;
      for (i = 1; i < 3; i = i + 1)
        s491 [i] <= s491 [i - 1];
      s493 [0] <= s795;
      for (i = 1; i < 3; i = i + 1)
        s493 [i] <= s493 [i - 1];
      s496 <= s761;
      s498 [0] <= s526;
      for (i = 1; i < 314; i = i + 1)
        s498 [i] <= s498 [i - 1];
      s499 <= s904;
      s500 <= s905;
      s504 [s186] <= s430;
      s503 <= s504 [s440];
      s506 [0] <= next;
      for (i = 1; i < 512; i = i + 1)
        s506 [i] <= s506 [i - 1];
      s507 <= s656;
      s509 [0] <= s884;
      for (i = 1; i < 15; i = i + 1)
        s509 [i] <= s509 [i - 1];
      s510 <= s781;
      s514 [0] <= s475;
      for (i = 1; i < 556; i = i + 1)
        s514 [i] <= s514 [i - 1];
      s515 <= s520;
      s517 [0] <= s358;
      for (i = 1; i < 3; i = i + 1)
        s517 [i] <= s517 [i - 1];
      s519 [0] <= s359;
      for (i = 1; i < 3; i = i + 1)
        s519 [i] <= s519 [i - 1];
      s522 [0] <= s346;
      for (i = 1; i < 10; i = i + 1)
        s522 [i] <= s522 [i - 1];
      s524 <= s193;
      s527 [0] <= s460;
      for (i = 1; i < 7; i = i + 1)
        s527 [i] <= s527 [i - 1];
      s529 [0] <= s615;
      for (i = 1; i < 12; i = i + 1)
        s529 [i] <= s529 [i - 1];
      s530 <= s260;
      s531 <= s944;
      s533 <= s32;
      s534 <= s731;
      s538 [0] <= s3;
      for (i = 1; i < 4; i = i + 1)
        s538 [i] <= s538 [i - 1];
      s540 <= s926;
      s542 [0] <= s472;
      for (i = 1; i < 518; i = i + 1)
        s542 [i] <= s542 [i - 1];
      s544 [0] <= s685;
      for (i = 1; i < 25; i = i + 1)
        s544 [i] <= s544 [i - 1];
      s545 <= s203;
      s547 [0] <= s533;
      for (i = 1; i < 127; i = i + 1)
        s547 [i] <= s547 [i - 1];
      s548 <= s426;
      s550 [0] <= s206;
      for (i = 1; i < 4; i = i + 1)
        s550 [i] <= s550 [i - 1];
      s553 <= s593;
      s555 [0] <= s248;
      for (i = 1; i < 4; i = i + 1)
        s555 [i] <= s555 [i - 1];
      s557 [0] <= s249;
      for (i = 1; i < 4; i = i + 1)
        s557 [i] <= s557 [i - 1];
      s559 <= s799;
      s558 <= s559;
      s561 <= s800;
      s560 <= s561;
      s566 [0] <= s417;
      for (i = 1; i < 255; i = i + 1)
        s566 [i] <= s566 [i - 1];
      s569 <= s582;
      s571 <= s933;
      s573 [0] <= s854;
      for (i = 1; i < 3; i = i + 1)
        s573 [i] <= s573 [i - 1];
      s575 [0] <= s855;
      for (i = 1; i < 3; i = i + 1)
        s575 [i] <= s575 [i - 1];
      s576 <= s299;
      s587 [0] <= s269;
      for (i = 1; i < 523; i = i + 1)
        s587 [i] <= s587 [i - 1];
      s589 <= s959;
      s588 <= s589;
      s591 <= s960;
      s590 <= s591;
      s595 [0] <= s850;
      for (i = 1; i < 265; i = i + 1)
        s595 [i] <= s595 [i - 1];
      s597 [0] <= s513;
      for (i = 1; i < 41; i = i + 1)
        s597 [i] <= s597 [i - 1];
      s606 <= s381;
      s607 <= s887;
      s609 <= s873;
      s610 <= s874;
      s612 [0] <= s327;
      for (i = 1; i < 6; i = i + 1)
        s612 [i] <= s612 [i - 1];
      s614 [0] <= s328;
      for (i = 1; i < 6; i = i + 1)
        s614 [i] <= s614 [i - 1];
      s616 [0] <= s726;
      for (i = 1; i < 17; i = i + 1)
        s616 [i] <= s616 [i - 1];
      s618 [0] <= s917;
      for (i = 1; i < 6; i = i + 1)
        s618 [i] <= s618 [i - 1];
      s622 <= s311;
      s623 <= s432;
      s624 <= s229;
      s625 <= s654;
      s627 [0] <= s35;
      for (i = 1; i < 4; i = i + 1)
        s627 [i] <= s627 [i - 1];
      s629 [0] <= s36;
      for (i = 1; i < 4; i = i + 1)
        s629 [i] <= s629 [i - 1];
      s633 [0] <= s48;
      for (i = 1; i < 132; i = i + 1)
        s633 [i] <= s633 [i - 1];
      s635 <= s892;
      s636 <= s893;
      s637 <= s747;
      s642 <= s211;
      s644 <= s176;
      s651 [0] <= s265;
      for (i = 1; i < 3; i = i + 1)
        s651 [i] <= s651 [i - 1];
      s653 [0] <= s266;
      for (i = 1; i < 3; i = i + 1)
        s653 [i] <= s653 [i - 1];
      s655 [s546] <= s5;
      s654 <= s655 [s533];
      s657 <= s797;
      s658 <= s953;
      s660 [0] <= s322;
      for (i = 1; i < 3; i = i + 1)
        s660 [i] <= s660 [i - 1];
      s662 [0] <= s323;
      for (i = 1; i < 3; i = i + 1)
        s662 [i] <= s662 [i - 1];
      s663 <= s108;
      s664 <= s109;
      s665 <= s495;
      s667 [0] <= s450;
      for (i = 1; i < 3; i = i + 1)
        s667 [i] <= s667 [i - 1];
      s669 [0] <= s451;
      for (i = 1; i < 3; i = i + 1)
        s669 [i] <= s669 [i - 1];
      s675 [0] <= s422;
      for (i = 1; i < 3; i = i + 1)
        s675 [i] <= s675 [i - 1];
      s677 [0] <= s423;
      for (i = 1; i < 3; i = i + 1)
        s677 [i] <= s677 [i - 1];
      s678 <= s836;
      s679 <= s293;
      s680 <= s230;
      s682 [0] <= s922;
      for (i = 1; i < 35; i = i + 1)
        s682 [i] <= s682 [i - 1];
      s683 <= s511;
      s684 <= s512;
      s686 [0] <= s476;
      for (i = 1; i < 546; i = i + 1)
        s686 [i] <= s686 [i - 1];
      s693 <= s945;
      s694 <= s579;
      s695 <= s580;
      s696 <= s640;
      s697 <= s641;
      s698 <= s635;
      s699 <= s636;
      s700 <= s885;
      s701 <= s307;
      s703 [0] <= s479;
      for (i = 1; i < 525; i = i + 1)
        s703 [i] <= s703 [i - 1];
      s704 <= s525;
      s711 [0] <= s43;
      for (i = 1; i < 4; i = i + 1)
        s711 [i] <= s711 [i - 1];
      s713 [0] <= s44;
      for (i = 1; i < 4; i = i + 1)
        s713 [i] <= s713 [i - 1];
      s715 <= s728;
      s719 [0] <= s254;
      for (i = 1; i < 63; i = i + 1)
        s719 [i] <= s719 [i - 1];
      s722 [0] <= s123;
      for (i = 1; i < 4; i = i + 1)
        s722 [i] <= s722 [i - 1];
      s724 [0] <= s124;
      for (i = 1; i < 4; i = i + 1)
        s724 [i] <= s724 [i - 1];
      s725 <= s409;
      s727 [0] <= s477;
      for (i = 1; i < 536; i = i + 1)
        s727 [i] <= s727 [i - 1];
      s730 [s279] <= s145;
      s729 <= s730 [s530];
      s732 <= s581;
      s738 [0] <= s235;
      for (i = 1; i < 63; i = i + 1)
        s738 [i] <= s738 [i - 1];
      s739 <= s37;
      s741 [0] <= s852;
      for (i = 1; i < 3; i = i + 1)
        s741 [i] <= s741 [i - 1];
      s743 [0] <= s853;
      for (i = 1; i < 3; i = i + 1)
        s743 [i] <= s743 [i - 1];
      s744 <= s437;
      s745 <= s1;
      s746 <= s2;
      s750 <= s687;
      s752 [0] <= s107;
      for (i = 1; i < 30; i = i + 1)
        s752 [i] <= s752 [i - 1];
      s753 <= s173;
      s754 <= s174;
      s756 <= s942;
      s757 <= s860;
      s758 <= s861;
      s759 <= s930;
      s760 <= s334;
      s763 [0] <= s715;
      for (i = 1; i < 7; i = i + 1)
        s763 [i] <= s763 [i - 1];
      s766 <= s568;
      s769 <= s643;
      s770 <= s362;
      s771 <= s363;
      s773 [0] <= s670;
      for (i = 1; i < 4; i = i + 1)
        s773 [i] <= s773 [i - 1];
      s775 [0] <= s671;
      for (i = 1; i < 4; i = i + 1)
        s775 [i] <= s775 [i - 1];
      s782 [0] <= s521;
      for (i = 1; i < 20; i = i + 1)
        s782 [i] <= s782 [i - 1];
      s784 [0] <= s645;
      for (i = 1; i < 3; i = i + 1)
        s784 [i] <= s784 [i - 1];
      s786 [0] <= s646;
      for (i = 1; i < 3; i = i + 1)
        s786 [i] <= s786 [i - 1];
      s788 [0] <= s324;
      for (i = 1; i < 4; i = i + 1)
        s788 [i] <= s788 [i - 1];
      s790 [0] <= s325;
      for (i = 1; i < 4; i = i + 1)
        s790 [i] <= s790 [i - 1];
      s796 <= s153;
      s799 <= s764;
      s800 <= s765;
      s801 <= s690;
      s803 [0] <= s318;
      for (i = 1; i < 250; i = i + 1)
        s803 [i] <= s803 [i - 1];
      s808 [0] <= s632;
      for (i = 1; i < 4; i = i + 1)
        s808 [i] <= s808 [i - 1];
      s814 <= s541;
      s813 <= s814;
      s819 <= s286;
      s818 <= s819;
      s821 <= s287;
      s820 <= s821;
      s823 [0] <= s200;
      for (i = 1; i < 4; i = i + 1)
        s823 [i] <= s823 [i - 1];
      s825 [0] <= s201;
      for (i = 1; i < 4; i = i + 1)
        s825 [i] <= s825 [i - 1];
      s826 <= s621;
      s827 <= s131;
      s830 <= s453;
      s831 <= s454;
      s832 <= s457;
      s834 <= s503;
      s838 [0] <= s76;
      for (i = 1; i < 16; i = i + 1)
        s838 [i] <= s838 [i - 1];
      s842 [0] <= s733;
      for (i = 1; i < 4; i = i + 1)
        s842 [i] <= s842 [i - 1];
      s844 [0] <= s734;
      for (i = 1; i < 4; i = i + 1)
        s844 [i] <= s844 [i - 1];
      s845 <= s644;
      s847 [0] <= s406;
      for (i = 1; i < 325; i = i + 1)
        s847 [i] <= s847 [i - 1];
      s851 [0] <= s902;
      for (i = 1; i < 70; i = i + 1)
        s851 [i] <= s851 [i - 1];
      s856 <= s197;
      s857 <= s867;
      s858 <= s868;
      s862 <= s501;
      s863 <= s502;
      s866 [0] <= s12;
      for (i = 1; i < 8; i = i + 1)
        s866 [i] <= s866 [i - 1];
      s869 <= s70;
      s871 [0] <= s596;
      for (i = 1; i < 36; i = i + 1)
        s871 [i] <= s871 [i - 1];
      s878 <= s111;
      s880 [0] <= s848;
      for (i = 1; i < 3; i = i + 1)
        s880 [i] <= s880 [i - 1];
      s882 [0] <= s849;
      for (i = 1; i < 3; i = i + 1)
        s882 [i] <= s882 [i - 1];
      s883 <= s16;
      s884 <= s243;
      s886 [s236] <= s170;
      s885 <= s886 [s606];
      s889 <= s270;
      s895 [0] <= s397;
      for (i = 1; i < 3; i = i + 1)
        s895 [i] <= s895 [i - 1];
      s897 [0] <= s398;
      for (i = 1; i < 3; i = i + 1)
        s897 [i] <= s897 [i - 1];
      s898 <= s805;
      s901 [0] <= s586;
      for (i = 1; i < 12; i = i + 1)
        s901 [i] <= s901 [i - 1];
      s903 [0] <= s22;
      for (i = 1; i < 485; i = i + 1)
        s903 [i] <= s903 [i - 1];
      s907 [0] <= s418;
      for (i = 1; i < 3; i = i + 1)
        s907 [i] <= s907 [i - 1];
      s910 <= s798;
      s914 <= s7;
      s916 [0] <= s681;
      for (i = 1; i < 228; i = i + 1)
        s916 [i] <= s916 [i - 1];
      s918 [0] <= s505;
      for (i = 1; i < 861; i = i + 1)
        s918 [i] <= s918 [i - 1];
      s923 [0] <= s524;
      for (i = 1; i < 31; i = i + 1)
        s923 [i] <= s923 [i - 1];
      s924 <= s345;
      s925 <= s673;
      s927 [s221] <= s68;
      s926 <= s927 [s239];
      s929 [0] <= s478;
      for (i = 1; i < 524; i = i + 1)
        s929 [i] <= s929 [i - 1];
      s932 [0] <= s305;
      for (i = 1; i < 154; i = i + 1)
        s932 [i] <= s932 [i - 1];
      s937 [0] <= s900;
      for (i = 1; i < 10; i = i + 1)
        s937 [i] <= s937 [i - 1];
      s938 <= s463;
      s940 [s288] <= s948;
      s939 <= s940 [s760];
      s943 [s737] <= s817;
      s942 <= s943 [s235];
      s947 [0] <= s845;
      for (i = 1; i < 338; i = i + 1)
        s947 [i] <= s947 [i - 1];
      s951 <= s872;
      s952 <= s608;
      s954 <= s238;
      s956 <= s857;
      s955 <= s956;
      s958 <= s858;
      s957 <= s958;
    end
endmodule

