module rgb_timing(
	input               i_rgb_clk,           //pixel clock
	input               i_rgb_rst_n,         //reset signal high active
	output  reg         o_rgb_hs,            //horizontal synchronization
	output  reg         o_rgb_vs,            //vertical synchronization
	output            	o_rgb_de,            //video valid

	output reg [10:0] 	o_rgb_x,              //video x position 
	output reg [10:0] 	o_rgb_y               //video y position 
	);


//800x480 33Mhz
parameter H_ACTIVE = 16'd800; 
parameter H_FP = 16'd40;      
parameter H_SYNC = 16'd128;   
parameter H_BP = 16'd88;      
parameter V_ACTIVE = 16'd480; 
parameter V_FP  = 16'd1;     
parameter V_SYNC  = 16'd3;    
parameter V_BP  = 16'd21;    
parameter HS_POL = 'b0;
parameter VS_POL = 'b0;

parameter H_TOTAL = H_ACTIVE + H_FP + H_SYNC + H_BP;//horizontal total time (pixels)
parameter V_TOTAL = V_ACTIVE + V_FP + V_SYNC + V_BP;//vertical total time (lines)

reg[11:0] h_cnt;                 //horizontal counter
reg[11:0] v_cnt;                 //vertical counter

reg h_active;                    //horizontal video active
reg v_active;                    //vertical video active
assign o_rgb_de = h_active & v_active;

always@(posedge i_rgb_clk)begin 
//显示计数
	if(h_cnt >= H_FP + H_SYNC + H_BP)
		o_rgb_x <= h_cnt - (H_FP[11:0] + H_SYNC[11:0] + H_BP[11:0]);
	else
		o_rgb_x <= o_rgb_x;
	if(v_cnt >= V_FP + V_SYNC + V_BP)
		o_rgb_y <= v_cnt - (V_FP[11:0] + V_SYNC[11:0] + V_BP[11:0]);
	else
		o_rgb_y <= o_rgb_y;
end

always@(posedge i_rgb_clk)begin 
//列计数
	if(i_rgb_rst_n == 'b0)
		h_cnt <= 'd0;
	else if(h_cnt == H_TOTAL - 1)//horizontal counter maximum value
		h_cnt <= 'd0;
	else
		h_cnt <= h_cnt + 'd1;
//行计数
	if(i_rgb_rst_n == 'b0)
		v_cnt <= 'd0;
	else if(h_cnt == H_FP  - 1)//horizontal sync time
		if(v_cnt == V_TOTAL - 1)//vertical counter maximum value
			v_cnt <= 'd0;
		else
			v_cnt <= v_cnt + 'd1;
	else
		v_cnt <= v_cnt;
//HS生成
	if(i_rgb_rst_n == 'b0)
		o_rgb_hs <= 'b0;
	else if(h_cnt == H_FP - 1)//horizontal sync begin
		o_rgb_hs <= HS_POL;
	else if(h_cnt == H_FP + H_SYNC - 1)//horizontal sync end
		o_rgb_hs <= ~o_rgb_hs;
	else
		o_rgb_hs <= o_rgb_hs;
//列有效
	if(i_rgb_rst_n == 'b0)
		h_active <= 'b0;
	else if(h_cnt == H_FP + H_SYNC + H_BP - 1)//horizontal active begin
		h_active <= 'b1;
	else if(h_cnt == H_TOTAL - 1)//horizontal active end
		h_active <= 'b0;
	else
		h_active <= h_active;
//VS生成
	if(i_rgb_rst_n == 'b0)
		o_rgb_vs <= 'd0;
	else if((v_cnt == V_FP - 1) && (h_cnt == H_FP - 1))//vertical sync begin
		o_rgb_vs <= VS_POL;
	else if((v_cnt == V_FP + V_SYNC - 1) && (h_cnt == H_FP - 1))//vertical sync end
		o_rgb_vs <= ~o_rgb_vs;  
	else
		o_rgb_vs <= o_rgb_vs;
//行有效
	if(i_rgb_rst_n == 'b0)
		v_active <= 'd0;
	else if((v_cnt == V_FP + V_SYNC + V_BP - 1) && (h_cnt == H_FP - 1))//vertical active begin
		v_active <= 'b1;
	else if((v_cnt == V_TOTAL - 1) && (h_cnt == H_FP - 1)) //vertical active end
		v_active <= 'b0;   
	else
		v_active <= v_active;
end
endmodule 