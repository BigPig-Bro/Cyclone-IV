module top(
    input           clk,

    output [9:0]    da5651e_db,
    output          da5651e_clk
);

parameter CLK_FRE 	= 50; //FPGA 输入MHz

/********************************************************************************/
/**************************      用户逻辑   ************************************/
/********************************************************************************/
wire [9:0] da5651e_data;
da5651e_ctl da5651e_ctl_m0(
    .clk            (clk            ),

    .da5651e_data   (da5651e_data    )
);

/********************************************************************************/
/**************************    da5651e驱动    ************************************/
/********************************************************************************/
assign da5651e_db    = da5651e_data;
assign da5651e_clk   = clk; //由于DAC clk频率通常较高，一般由PLL单独给出

endmodule